-- 32 Kbyte Block RAM, one R/W port, one read-only port

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity VideoRam is
generic (
	ADDR_BITS		: integer := 15;
	DATA_BITS		: integer := 8
);
port (
	Clock			: in  std_logic;
	Enable			: in  std_logic;
	WriteEnable		: in  std_logic;
	Address			: in  std_logic_vector(ADDR_BITS-1 downto 0);
	DataIn			: in  std_logic_vector(DATA_BITS-1 downto 0);
	DataOut			: out std_logic_vector(DATA_BITS-1 downto 0);

	DualEnable		: in  std_logic;
	DualAddress		: in  std_logic_vector(ADDR_BITS-1 downto 0);
	DualDataOut		: out std_logic_vector(DATA_BITS-1 downto 0)
);
end VideoRam;

architecture behavioral of VideoRam is

type ram_type is array (0 to 2**ADDR_BITS - 1) of std_logic_vector (DataOut'range);
signal RAM: ram_type := (

	x"f3",x"31",x"00",x"5c",x"af",x"d3",x"1f",x"3e",x"01",x"d3",x"fe",x"cd",x"f1",x"00",x"3a",x"25",
	x"05",x"fe",x"01",x"28",x"1c",x"3e",x"02",x"d3",x"fe",x"21",x"26",x"05",x"11",x"00",x"80",x"01",
	x"00",x"40",x"ed",x"b0",x"21",x"26",x"05",x"01",x"00",x"40",x"ed",x"b0",x"3e",x"01",x"32",x"25",
	x"05",x"21",x"00",x"40",x"22",x"00",x"5b",x"11",x"01",x"40",x"01",x"00",x"18",x"af",x"77",x"ed",
	x"b0",x"01",x"00",x"02",x"3e",x"78",x"77",x"ed",x"b0",x"06",x"40",x"af",x"77",x"23",x"77",x"23",
	x"77",x"23",x"77",x"23",x"c6",x"08",x"e6",x"7f",x"10",x"f2",x"11",x"61",x"04",x"cd",x"21",x"01",
	x"01",x"c8",x"00",x"2e",x"07",x"7d",x"d3",x"fe",x"ee",x"10",x"6f",x"c5",x"06",x"64",x"10",x"fe",
	x"c1",x"0b",x"78",x"b1",x"20",x"ef",x"01",x"fe",x"f7",x"ed",x"78",x"2f",x"e6",x"1f",x"32",x"02",
	x"5b",x"b7",x"28",x"f2",x"ed",x"78",x"e6",x"1f",x"fe",x"1f",x"20",x"f8",x"3a",x"02",x"5b",x"fe",
	x"10",x"28",x"1a",x"fe",x"01",x"26",x"00",x"28",x"20",x"fe",x"02",x"26",x"40",x"28",x"1a",x"fe",
	x"04",x"26",x"80",x"28",x"14",x"fe",x"08",x"26",x"c0",x"28",x"0e",x"18",x"c9",x"11",x"05",x"05",
	x"cd",x"21",x"01",x"3e",x"03",x"d3",x"fe",x"18",x"44",x"11",x"12",x"05",x"cd",x"21",x"01",x"3e",
	x"04",x"d3",x"fe",x"3e",x"03",x"d3",x"1f",x"3e",x"03",x"d3",x"3f",x"3e",x"3f",x"d3",x"3f",x"7c",
	x"d3",x"3f",x"af",x"d3",x"3f",x"01",x"00",x"80",x"11",x"00",x"80",x"d3",x"3f",x"db",x"3f",x"12",
	x"13",x"0b",x"78",x"b1",x"20",x"f5",x"af",x"d3",x"1f",x"11",x"20",x"05",x"cd",x"21",x"01",x"18",
	x"0c",x"01",x"fd",x"42",x"3e",x"80",x"ed",x"79",x"3e",x"c1",x"ed",x"79",x"c9",x"21",x"0b",x"01",
	x"11",x"00",x"5c",x"01",x"16",x"00",x"ed",x"b0",x"c3",x"00",x"5c",x"3e",x"06",x"d3",x"fe",x"01",
	x"fd",x"42",x"3e",x"20",x"ed",x"79",x"3e",x"82",x"ed",x"79",x"3e",x"c3",x"ed",x"79",x"c3",x"00",
	x"00",x"1a",x"b7",x"c8",x"13",x"cd",x"2a",x"01",x"18",x"f7",x"d9",x"fe",x"0a",x"28",x"1e",x"6f",
	x"26",x"00",x"29",x"29",x"29",x"11",x"61",x"00",x"19",x"ed",x"5b",x"00",x"5b",x"13",x"ed",x"53",
	x"00",x"5b",x"1b",x"06",x"08",x"7e",x"12",x"23",x"14",x"10",x"fa",x"18",x"12",x"2a",x"00",x"5b",
	x"7d",x"e6",x"e0",x"c6",x"20",x"6f",x"30",x"04",x"7c",x"c6",x"08",x"67",x"22",x"00",x"5b",x"d9",
	x"c9",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"00",x"10",
	x"00",x"00",x"6c",x"24",x"48",x"00",x"00",x"00",x"00",x"00",x"28",x"7c",x"28",x"28",x"7c",x"28",
	x"00",x"00",x"10",x"3c",x"40",x"38",x"04",x"78",x"10",x"00",x"42",x"a4",x"48",x"10",x"24",x"4a",
	x"84",x"00",x"30",x"40",x"36",x"44",x"44",x"38",x"00",x"00",x"18",x"08",x"10",x"00",x"00",x"00",
	x"00",x"00",x"08",x"10",x"10",x"10",x"10",x"10",x"08",x"00",x"20",x"10",x"10",x"10",x"10",x"10",
	x"20",x"00",x"00",x"28",x"10",x"7c",x"10",x"28",x"00",x"00",x"00",x"10",x"10",x"7c",x"10",x"10",
	x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"08",x"10",x"00",x"00",x"00",x"00",x"7c",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"00",x"00",x"02",x"04",x"08",x"10",x"20",x"40",
	x"00",x"00",x"38",x"44",x"54",x"54",x"44",x"38",x"00",x"00",x"10",x"70",x"10",x"10",x"10",x"7c",
	x"00",x"00",x"38",x"44",x"04",x"38",x"40",x"7c",x"00",x"00",x"38",x"44",x"18",x"04",x"44",x"38",
	x"00",x"00",x"18",x"28",x"28",x"48",x"7c",x"08",x"00",x"00",x"7c",x"40",x"78",x"04",x"44",x"38",
	x"00",x"00",x"38",x"40",x"78",x"44",x"44",x"38",x"00",x"00",x"7c",x"04",x"08",x"08",x"10",x"10",
	x"00",x"00",x"38",x"44",x"38",x"44",x"44",x"38",x"00",x"00",x"38",x"44",x"44",x"3c",x"04",x"38",
	x"00",x"00",x"00",x"10",x"10",x"00",x"10",x"10",x"00",x"00",x"00",x"10",x"10",x"00",x"30",x"10",
	x"20",x"00",x"00",x"08",x"10",x"20",x"10",x"08",x"00",x"00",x"00",x"00",x"7c",x"00",x"7c",x"00",
	x"00",x"00",x"00",x"10",x"08",x"04",x"08",x"10",x"00",x"00",x"38",x"04",x"08",x"10",x"00",x"10",
	x"00",x"00",x"38",x"44",x"92",x"aa",x"9c",x"40",x"3c",x"00",x"38",x"44",x"44",x"7c",x"44",x"44",
	x"00",x"00",x"78",x"44",x"78",x"44",x"44",x"78",x"00",x"00",x"38",x"44",x"40",x"40",x"44",x"38",
	x"00",x"00",x"78",x"44",x"44",x"44",x"44",x"78",x"00",x"00",x"3c",x"20",x"3c",x"20",x"20",x"3c",
	x"00",x"00",x"3c",x"20",x"20",x"3c",x"20",x"20",x"00",x"00",x"38",x"44",x"40",x"4c",x"44",x"3c",
	x"00",x"00",x"44",x"44",x"7c",x"44",x"44",x"44",x"00",x"00",x"38",x"10",x"10",x"10",x"10",x"38",
	x"00",x"00",x"04",x"04",x"04",x"44",x"44",x"38",x"00",x"00",x"44",x"48",x"50",x"70",x"48",x"44",
	x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"3c",x"00",x"00",x"44",x"6c",x"54",x"44",x"44",x"44",
	x"00",x"00",x"44",x"64",x"54",x"4c",x"44",x"44",x"00",x"00",x"38",x"44",x"44",x"44",x"44",x"38",
	x"00",x"00",x"78",x"44",x"44",x"58",x"40",x"40",x"00",x"00",x"38",x"44",x"44",x"44",x"44",x"38",
	x"04",x"00",x"78",x"44",x"44",x"78",x"48",x"44",x"00",x"00",x"38",x"40",x"38",x"04",x"44",x"38",
	x"00",x"00",x"7c",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"44",x"44",x"44",x"44",x"44",x"38",
	x"00",x"00",x"44",x"44",x"28",x"28",x"10",x"10",x"00",x"00",x"44",x"44",x"54",x"54",x"54",x"28",
	x"00",x"00",x"44",x"28",x"10",x"10",x"28",x"44",x"00",x"00",x"44",x"44",x"28",x"10",x"10",x"10",
	x"00",x"00",x"3c",x"04",x"08",x"10",x"20",x"3c",x"00",x"00",x"18",x"10",x"10",x"10",x"10",x"10",
	x"18",x"00",x"40",x"20",x"10",x"08",x"04",x"02",x"00",x"00",x"30",x"10",x"10",x"10",x"10",x"10",
	x"30",x"00",x"10",x"28",x"44",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"7e",x"00",x"18",x"20",x"78",x"20",x"20",x"7c",x"00",x"00",x"00",x"38",x"04",x"3c",x"44",x"3c",
	x"00",x"00",x"40",x"58",x"64",x"44",x"44",x"78",x"00",x"00",x"00",x"38",x"40",x"40",x"44",x"38",
	x"00",x"00",x"04",x"34",x"4c",x"44",x"44",x"3c",x"00",x"00",x"00",x"38",x"44",x"7c",x"40",x"38",
	x"00",x"00",x"0c",x"10",x"7c",x"10",x"10",x"10",x"00",x"00",x"00",x"3c",x"44",x"4c",x"34",x"04",
	x"38",x"00",x"40",x"58",x"64",x"44",x"44",x"44",x"00",x"00",x"10",x"00",x"70",x"10",x"10",x"10",
	x"00",x"00",x"08",x"00",x"38",x"08",x"08",x"08",x"70",x"00",x"40",x"44",x"48",x"70",x"48",x"44",
	x"00",x"00",x"20",x"20",x"20",x"20",x"24",x"18",x"00",x"00",x"00",x"ec",x"92",x"92",x"92",x"92",
	x"00",x"00",x"00",x"58",x"64",x"44",x"44",x"44",x"00",x"00",x"00",x"38",x"44",x"44",x"44",x"38",
	x"00",x"00",x"00",x"58",x"64",x"44",x"44",x"78",x"40",x"00",x"00",x"3c",x"44",x"44",x"4c",x"34",
	x"04",x"00",x"00",x"2c",x"30",x"20",x"20",x"20",x"00",x"00",x"00",x"38",x"40",x"38",x"04",x"78",
	x"00",x"00",x"20",x"7c",x"20",x"20",x"24",x"18",x"00",x"00",x"00",x"44",x"44",x"44",x"4c",x"34",
	x"00",x"00",x"00",x"44",x"44",x"28",x"28",x"10",x"00",x"00",x"00",x"92",x"92",x"92",x"92",x"6c",
	x"00",x"00",x"00",x"44",x"28",x"10",x"28",x"44",x"00",x"00",x"00",x"44",x"44",x"28",x"28",x"10",
	x"60",x"00",x"00",x"7c",x"08",x"10",x"20",x"7c",x"00",x"00",x"08",x"10",x"10",x"20",x"10",x"10",
	x"08",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"20",x"10",x"10",x"08",x"10",x"10",
	x"20",x"00",x"34",x"58",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"44",x"92",x"a2",x"92",x"44",
	x"38",x"48",x"43",x"2d",x"46",x"6f",x"72",x"65",x"76",x"65",x"72",x"20",x"28",x"72",x"65",x"76",
	x"20",x"42",x"29",x"0a",x"43",x"6f",x"70",x"79",x"72",x"69",x"67",x"68",x"74",x"20",x"7f",x"20",
	x"32",x"30",x"30",x"35",x"2d",x"32",x"30",x"31",x"32",x"20",x"41",x"6c",x"65",x"78",x"20",x"42",
	x"61",x"64",x"65",x"61",x"20",x"3c",x"76",x"61",x"6d",x"70",x"6f",x"73",x"64",x"65",x"63",x"61",
	x"6d",x"70",x"6f",x"73",x"40",x"67",x"6d",x"61",x"69",x"6c",x"2e",x"63",x"6f",x"6d",x"3e",x"0a",
	x"0a",x"42",x"6f",x"6f",x"74",x"6c",x"6f",x"61",x"64",x"65",x"72",x"20",x"34",x"33",x"63",x"37",
	x"30",x"39",x"65",x"33",x"20",x"2f",x"20",x"32",x"30",x"31",x"32",x"2d",x"30",x"32",x"2d",x"32",
	x"33",x"43",x"68",x"6f",x"6f",x"73",x"65",x"20",x"69",x"6d",x"61",x"67",x"65",x"3a",x"0a",x"20",
	x"20",x"31",x"2e",x"2e",x"34",x"20",x"2d",x"20",x"53",x"50",x"49",x"20",x"66",x"6c",x"61",x"73",
	x"68",x"0a",x"20",x"20",x"35",x"20",x"20",x"20",x"20",x"2d",x"20",x"6d",x"61",x"73",x"6b",x"20",
	x"52",x"4f",x"4d",x"0a",x"00",x"6d",x"61",x"73",x"6b",x"20",x"52",x"4f",x"4d",x"2e",x"2e",x"2e",
	x"20",x"00",x"53",x"50",x"49",x"20",x"66",x"6c",x"61",x"73",x"68",x"2e",x"2e",x"2e",x"20",x"00",
	x"64",x"6f",x"6e",x"65",x"00",x"00",x"f3",x"af",x"11",x"ff",x"ff",x"c3",x"cb",x"11",x"2a",x"5d",
	x"5c",x"22",x"5f",x"5c",x"18",x"43",x"c3",x"f2",x"15",x"ff",x"ff",x"ff",x"ff",x"ff",x"2a",x"5d",
	x"5c",x"7e",x"cd",x"7d",x"00",x"d0",x"cd",x"74",x"00",x"18",x"f7",x"ff",x"ff",x"ff",x"c3",x"5b",
	x"33",x"ff",x"ff",x"ff",x"ff",x"ff",x"c5",x"2a",x"61",x"5c",x"e5",x"c3",x"9e",x"16",x"f5",x"e5",
	x"2a",x"78",x"5c",x"23",x"22",x"78",x"5c",x"7c",x"b5",x"20",x"03",x"fd",x"34",x"40",x"c5",x"d5",
	x"cd",x"bf",x"02",x"d1",x"c1",x"e1",x"f1",x"fb",x"c9",x"e1",x"6e",x"fd",x"75",x"00",x"ed",x"7b",
	x"3d",x"5c",x"c3",x"c5",x"16",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f5",x"e5",x"2a",x"b0",
	x"5c",x"7c",x"b5",x"20",x"01",x"e9",x"e1",x"f1",x"ed",x"45",x"2a",x"5d",x"5c",x"23",x"22",x"5d",
	x"5c",x"7e",x"c9",x"fe",x"21",x"d0",x"fe",x"0d",x"c8",x"fe",x"10",x"d8",x"fe",x"18",x"3f",x"d8",
	x"23",x"fe",x"16",x"38",x"01",x"23",x"37",x"22",x"5d",x"5c",x"c9",x"bf",x"52",x"4e",x"c4",x"49",
	x"4e",x"4b",x"45",x"59",x"a4",x"50",x"c9",x"46",x"ce",x"50",x"4f",x"49",x"4e",x"d4",x"53",x"43",
	x"52",x"45",x"45",x"4e",x"a4",x"41",x"54",x"54",x"d2",x"41",x"d4",x"54",x"41",x"c2",x"56",x"41",
	x"4c",x"a4",x"43",x"4f",x"44",x"c5",x"56",x"41",x"cc",x"4c",x"45",x"ce",x"53",x"49",x"ce",x"43",
	x"4f",x"d3",x"54",x"41",x"ce",x"41",x"53",x"ce",x"41",x"43",x"d3",x"41",x"54",x"ce",x"4c",x"ce",
	x"45",x"58",x"d0",x"49",x"4e",x"d4",x"53",x"51",x"d2",x"53",x"47",x"ce",x"41",x"42",x"d3",x"50",
	x"45",x"45",x"cb",x"49",x"ce",x"55",x"53",x"d2",x"53",x"54",x"52",x"a4",x"43",x"48",x"52",x"a4",
	x"4e",x"4f",x"d4",x"42",x"49",x"ce",x"4f",x"d2",x"41",x"4e",x"c4",x"3c",x"bd",x"3e",x"bd",x"3c",
	x"be",x"4c",x"49",x"4e",x"c5",x"54",x"48",x"45",x"ce",x"54",x"cf",x"53",x"54",x"45",x"d0",x"44",
	x"45",x"46",x"20",x"46",x"ce",x"43",x"41",x"d4",x"46",x"4f",x"52",x"4d",x"41",x"d4",x"4d",x"4f",
	x"56",x"c5",x"45",x"52",x"41",x"53",x"c5",x"4f",x"50",x"45",x"4e",x"20",x"a3",x"43",x"4c",x"4f",
	x"53",x"45",x"20",x"a3",x"4d",x"45",x"52",x"47",x"c5",x"56",x"45",x"52",x"49",x"46",x"d9",x"42",
	x"45",x"45",x"d0",x"43",x"49",x"52",x"43",x"4c",x"c5",x"49",x"4e",x"cb",x"50",x"41",x"50",x"45",
	x"d2",x"46",x"4c",x"41",x"53",x"c8",x"42",x"52",x"49",x"47",x"48",x"d4",x"49",x"4e",x"56",x"45",
	x"52",x"53",x"c5",x"4f",x"56",x"45",x"d2",x"4f",x"55",x"d4",x"4c",x"50",x"52",x"49",x"4e",x"d4",
	x"4c",x"4c",x"49",x"53",x"d4",x"53",x"54",x"4f",x"d0",x"52",x"45",x"41",x"c4",x"44",x"41",x"54",
	x"c1",x"52",x"45",x"53",x"54",x"4f",x"52",x"c5",x"4e",x"45",x"d7",x"42",x"4f",x"52",x"44",x"45",
	x"d2",x"43",x"4f",x"4e",x"54",x"49",x"4e",x"55",x"c5",x"44",x"49",x"cd",x"52",x"45",x"cd",x"46",
	x"4f",x"d2",x"47",x"4f",x"20",x"54",x"cf",x"47",x"4f",x"20",x"53",x"55",x"c2",x"49",x"4e",x"50",
	x"55",x"d4",x"4c",x"4f",x"41",x"c4",x"4c",x"49",x"53",x"d4",x"4c",x"45",x"d4",x"50",x"41",x"55",
	x"53",x"c5",x"4e",x"45",x"58",x"d4",x"50",x"4f",x"4b",x"c5",x"50",x"52",x"49",x"4e",x"d4",x"50",
	x"4c",x"4f",x"d4",x"52",x"55",x"ce",x"53",x"41",x"56",x"c5",x"52",x"41",x"4e",x"44",x"4f",x"4d",
	x"49",x"5a",x"c5",x"49",x"c6",x"43",x"4c",x"d3",x"44",x"52",x"41",x"d7",x"43",x"4c",x"45",x"41",
	x"d2",x"52",x"45",x"54",x"55",x"52",x"ce",x"43",x"4f",x"50",x"d9",x"42",x"48",x"59",x"36",x"35",
	x"54",x"47",x"56",x"4e",x"4a",x"55",x"37",x"34",x"52",x"46",x"43",x"4d",x"4b",x"49",x"38",x"33",
	x"45",x"44",x"58",x"0e",x"4c",x"4f",x"39",x"32",x"57",x"53",x"5a",x"20",x"0d",x"50",x"30",x"31",
	x"51",x"41",x"e3",x"c4",x"e0",x"e4",x"b4",x"bc",x"bd",x"bb",x"af",x"b0",x"b1",x"c0",x"a7",x"a6",
	x"be",x"ad",x"b2",x"ba",x"e5",x"a5",x"c2",x"e1",x"b3",x"b9",x"c1",x"b8",x"7e",x"dc",x"da",x"5c",
	x"b7",x"7b",x"7d",x"d8",x"bf",x"ae",x"aa",x"ab",x"dd",x"de",x"df",x"7f",x"b5",x"d6",x"7c",x"d5",
	x"5d",x"db",x"b6",x"d9",x"5b",x"d7",x"0c",x"07",x"06",x"04",x"05",x"08",x"0a",x"0b",x"09",x"0f",
	x"e2",x"2a",x"3f",x"cd",x"c8",x"cc",x"cb",x"5e",x"ac",x"2d",x"2b",x"3d",x"2e",x"2c",x"3b",x"22",
	x"c7",x"3c",x"c3",x"3e",x"c5",x"2f",x"c9",x"60",x"c6",x"3a",x"d0",x"ce",x"a8",x"ca",x"d3",x"d4",
	x"d1",x"d2",x"a9",x"cf",x"2e",x"2f",x"11",x"ff",x"ff",x"01",x"fe",x"fe",x"ed",x"78",x"2f",x"e6",
	x"1f",x"28",x"0e",x"67",x"7d",x"14",x"c0",x"d6",x"08",x"cb",x"3c",x"30",x"fa",x"53",x"5f",x"20",
	x"f4",x"2d",x"cb",x"00",x"38",x"e6",x"7a",x"3c",x"c8",x"fe",x"28",x"c8",x"fe",x"19",x"c8",x"7b",
	x"5a",x"57",x"fe",x"18",x"c9",x"cd",x"8e",x"02",x"c0",x"21",x"00",x"5c",x"cb",x"7e",x"20",x"07",
	x"23",x"35",x"2b",x"20",x"02",x"36",x"ff",x"7d",x"21",x"04",x"5c",x"bd",x"20",x"ee",x"cd",x"1e",
	x"03",x"d0",x"21",x"00",x"5c",x"be",x"28",x"2e",x"eb",x"21",x"04",x"5c",x"be",x"28",x"27",x"cb",
	x"7e",x"20",x"04",x"eb",x"cb",x"7e",x"c8",x"5f",x"77",x"23",x"36",x"05",x"23",x"3a",x"09",x"5c",
	x"77",x"23",x"fd",x"4e",x"07",x"fd",x"56",x"01",x"e5",x"cd",x"33",x"03",x"e1",x"77",x"32",x"08",
	x"5c",x"fd",x"cb",x"01",x"ee",x"c9",x"23",x"36",x"05",x"23",x"35",x"c0",x"3a",x"0a",x"5c",x"77",
	x"23",x"7e",x"18",x"ea",x"42",x"16",x"00",x"7b",x"fe",x"27",x"d0",x"fe",x"18",x"20",x"03",x"cb",
	x"78",x"c0",x"21",x"05",x"02",x"19",x"7e",x"37",x"c9",x"7b",x"fe",x"3a",x"38",x"2f",x"0d",x"fa",
	x"4f",x"03",x"28",x"03",x"c6",x"4f",x"c9",x"21",x"eb",x"01",x"04",x"28",x"03",x"21",x"05",x"02",
	x"16",x"00",x"19",x"7e",x"c9",x"21",x"29",x"02",x"cb",x"40",x"28",x"f4",x"cb",x"5a",x"28",x"0a",
	x"fd",x"cb",x"30",x"5e",x"c0",x"04",x"c0",x"c6",x"20",x"c9",x"c6",x"a5",x"c9",x"fe",x"30",x"d8",
	x"0d",x"fa",x"9d",x"03",x"20",x"19",x"21",x"54",x"02",x"cb",x"68",x"28",x"d3",x"fe",x"38",x"30",
	x"07",x"d6",x"20",x"04",x"c8",x"c6",x"08",x"c9",x"d6",x"36",x"04",x"c8",x"c6",x"fe",x"c9",x"21",
	x"30",x"02",x"fe",x"39",x"28",x"ba",x"fe",x"30",x"28",x"b6",x"e6",x"07",x"c6",x"80",x"04",x"c8",
	x"ee",x"0f",x"c9",x"04",x"c8",x"cb",x"68",x"21",x"30",x"02",x"20",x"a4",x"d6",x"10",x"fe",x"22",
	x"28",x"06",x"fe",x"20",x"c0",x"3e",x"5f",x"c9",x"3e",x"40",x"c9",x"f3",x"7d",x"cb",x"3d",x"cb",
	x"3d",x"2f",x"e6",x"03",x"4f",x"06",x"00",x"dd",x"21",x"d1",x"03",x"dd",x"09",x"3a",x"48",x"5c",
	x"e6",x"38",x"0f",x"0f",x"0f",x"f6",x"08",x"00",x"00",x"00",x"04",x"0c",x"0d",x"20",x"fd",x"0e",
	x"3f",x"05",x"c2",x"d6",x"03",x"ee",x"10",x"d3",x"fe",x"44",x"4f",x"cb",x"67",x"20",x"09",x"7a",
	x"b3",x"28",x"09",x"79",x"4d",x"1b",x"dd",x"e9",x"4d",x"0c",x"dd",x"e9",x"fb",x"c9",x"ef",x"31",
	x"27",x"c0",x"03",x"34",x"ec",x"6c",x"98",x"1f",x"f5",x"04",x"a1",x"0f",x"38",x"21",x"92",x"5c",
	x"7e",x"a7",x"20",x"5e",x"23",x"4e",x"23",x"46",x"78",x"17",x"9f",x"b9",x"20",x"54",x"23",x"be",
	x"20",x"50",x"78",x"c6",x"3c",x"f2",x"25",x"04",x"e2",x"6c",x"04",x"06",x"fa",x"04",x"d6",x"0c",
	x"30",x"fb",x"c6",x"0c",x"c5",x"21",x"6e",x"04",x"cd",x"06",x"34",x"cd",x"b4",x"33",x"ef",x"04",
	x"38",x"f1",x"86",x"77",x"ef",x"c0",x"02",x"31",x"38",x"cd",x"94",x"1e",x"fe",x"0b",x"30",x"22",
	x"ef",x"e0",x"04",x"e0",x"34",x"80",x"43",x"55",x"9f",x"80",x"01",x"05",x"34",x"35",x"71",x"03",
	x"38",x"cd",x"99",x"1e",x"c5",x"cd",x"99",x"1e",x"e1",x"50",x"59",x"7a",x"b3",x"c8",x"1b",x"c3",
	x"b5",x"03",x"cf",x"0a",x"89",x"02",x"d0",x"12",x"86",x"89",x"0a",x"97",x"60",x"75",x"89",x"12",
	x"d5",x"17",x"1f",x"89",x"1b",x"90",x"41",x"02",x"89",x"24",x"d0",x"53",x"ca",x"89",x"2e",x"9d",
	x"36",x"b1",x"89",x"38",x"ff",x"49",x"3e",x"89",x"43",x"ff",x"6a",x"73",x"89",x"4f",x"a7",x"00",
	x"54",x"89",x"5c",x"00",x"00",x"00",x"89",x"69",x"14",x"f6",x"24",x"89",x"76",x"f1",x"10",x"05",
	x"cd",x"fb",x"24",x"3a",x"3b",x"5c",x"87",x"fa",x"8a",x"1c",x"e1",x"d0",x"e5",x"cd",x"f1",x"2b",
	x"62",x"6b",x"0d",x"f8",x"09",x"cb",x"fe",x"c9",x"21",x"3f",x"05",x"e5",x"21",x"80",x"1f",x"cb",
	x"7f",x"28",x"03",x"21",x"98",x"0c",x"08",x"13",x"dd",x"2b",x"f3",x"3e",x"02",x"47",x"10",x"fe",
	x"d3",x"fe",x"ee",x"0f",x"06",x"a4",x"2d",x"20",x"f5",x"05",x"25",x"f2",x"d8",x"04",x"06",x"2f",
	x"10",x"fe",x"d3",x"fe",x"3e",x"0d",x"06",x"37",x"10",x"fe",x"d3",x"fe",x"01",x"0e",x"3b",x"08",
	x"6f",x"c3",x"07",x"05",x"7a",x"b3",x"28",x"0c",x"dd",x"6e",x"00",x"7c",x"ad",x"67",x"3e",x"01",
	x"37",x"c3",x"25",x"05",x"6c",x"18",x"f4",x"79",x"cb",x"78",x"10",x"fe",x"30",x"04",x"06",x"42",
	x"10",x"fe",x"d3",x"fe",x"06",x"3e",x"20",x"ef",x"05",x"af",x"3c",x"cb",x"15",x"c2",x"14",x"05",
	x"1b",x"dd",x"23",x"06",x"31",x"3e",x"7f",x"db",x"fe",x"1f",x"d0",x"7a",x"3c",x"c2",x"fe",x"04",
	x"06",x"3b",x"10",x"fe",x"c9",x"f5",x"3a",x"48",x"5c",x"e6",x"38",x"0f",x"0f",x"0f",x"d3",x"fe",
	x"3e",x"7f",x"db",x"fe",x"1f",x"fb",x"38",x"02",x"cf",x"0c",x"f1",x"c9",x"14",x"08",x"15",x"f3",
	x"3e",x"0f",x"d3",x"fe",x"21",x"3f",x"05",x"e5",x"db",x"fe",x"1f",x"e6",x"20",x"f6",x"02",x"4f",
	x"bf",x"c0",x"cd",x"e7",x"05",x"30",x"fa",x"21",x"15",x"04",x"10",x"fe",x"2b",x"7c",x"b5",x"20",
	x"f9",x"cd",x"e3",x"05",x"30",x"eb",x"06",x"9c",x"cd",x"e3",x"05",x"30",x"e4",x"3e",x"c6",x"b8",
	x"30",x"e0",x"24",x"20",x"f1",x"06",x"c9",x"cd",x"e7",x"05",x"30",x"d5",x"78",x"fe",x"d4",x"30",
	x"f4",x"cd",x"e7",x"05",x"d0",x"79",x"ee",x"03",x"4f",x"26",x"00",x"06",x"b0",x"18",x"1f",x"08",
	x"20",x"07",x"30",x"0f",x"dd",x"75",x"00",x"18",x"0f",x"cb",x"11",x"ad",x"c0",x"79",x"1f",x"4f",
	x"13",x"18",x"07",x"dd",x"7e",x"00",x"ad",x"c0",x"dd",x"23",x"1b",x"08",x"06",x"b2",x"2e",x"01",
	x"cd",x"e3",x"05",x"d0",x"3e",x"cb",x"b8",x"cb",x"15",x"06",x"b0",x"d2",x"ca",x"05",x"7c",x"ad",
	x"67",x"7a",x"b3",x"20",x"ca",x"7c",x"fe",x"01",x"c9",x"cd",x"e7",x"05",x"d0",x"3e",x"16",x"3d",
	x"20",x"fd",x"a7",x"04",x"c8",x"3e",x"7f",x"db",x"fe",x"1f",x"d0",x"a9",x"e6",x"20",x"28",x"f3",
	x"79",x"2f",x"4f",x"e6",x"07",x"f6",x"08",x"d3",x"fe",x"37",x"c9",x"f1",x"3a",x"74",x"5c",x"d6",
	x"e0",x"32",x"74",x"5c",x"cd",x"8c",x"1c",x"cd",x"30",x"25",x"28",x"3c",x"01",x"11",x"00",x"3a",
	x"74",x"5c",x"a7",x"28",x"02",x"0e",x"22",x"f7",x"d5",x"dd",x"e1",x"06",x"0b",x"3e",x"20",x"12",
	x"13",x"10",x"fc",x"dd",x"36",x"01",x"ff",x"cd",x"f1",x"2b",x"21",x"f6",x"ff",x"0b",x"09",x"03",
	x"30",x"0f",x"3a",x"74",x"5c",x"a7",x"20",x"02",x"cf",x"0e",x"78",x"b1",x"28",x"0a",x"01",x"0a",
	x"00",x"dd",x"e5",x"e1",x"23",x"eb",x"ed",x"b0",x"df",x"fe",x"e4",x"20",x"49",x"3a",x"74",x"5c",
	x"fe",x"03",x"ca",x"8a",x"1c",x"e7",x"cd",x"b2",x"28",x"cb",x"f9",x"30",x"0b",x"21",x"00",x"00",
	x"3a",x"74",x"5c",x"3d",x"28",x"15",x"cf",x"01",x"c2",x"8a",x"1c",x"cd",x"30",x"25",x"28",x"18",
	x"23",x"7e",x"dd",x"77",x"0b",x"23",x"7e",x"dd",x"77",x"0c",x"23",x"dd",x"71",x"0e",x"3e",x"01",
	x"cb",x"71",x"28",x"01",x"3c",x"dd",x"77",x"00",x"eb",x"e7",x"fe",x"29",x"20",x"da",x"e7",x"cd",
	x"ee",x"1b",x"eb",x"c3",x"5a",x"07",x"fe",x"aa",x"20",x"1f",x"3a",x"74",x"5c",x"fe",x"03",x"ca",
	x"8a",x"1c",x"e7",x"cd",x"ee",x"1b",x"dd",x"36",x"0b",x"00",x"dd",x"36",x"0c",x"1b",x"21",x"00",
	x"40",x"dd",x"75",x"0d",x"dd",x"74",x"0e",x"18",x"4d",x"fe",x"af",x"20",x"4f",x"3a",x"74",x"5c",
	x"fe",x"03",x"ca",x"8a",x"1c",x"e7",x"cd",x"48",x"20",x"20",x"0c",x"3a",x"74",x"5c",x"a7",x"ca",
	x"8a",x"1c",x"cd",x"e6",x"1c",x"18",x"0f",x"cd",x"82",x"1c",x"df",x"fe",x"2c",x"28",x"0c",x"3a",
	x"74",x"5c",x"a7",x"ca",x"8a",x"1c",x"cd",x"e6",x"1c",x"18",x"04",x"e7",x"cd",x"82",x"1c",x"cd",
	x"ee",x"1b",x"cd",x"99",x"1e",x"dd",x"71",x"0b",x"dd",x"70",x"0c",x"cd",x"99",x"1e",x"dd",x"71",
	x"0d",x"dd",x"70",x"0e",x"60",x"69",x"dd",x"36",x"00",x"03",x"18",x"44",x"fe",x"ca",x"28",x"09",
	x"cd",x"ee",x"1b",x"dd",x"36",x"0e",x"80",x"18",x"17",x"3a",x"74",x"5c",x"a7",x"c2",x"8a",x"1c",
	x"e7",x"cd",x"82",x"1c",x"cd",x"ee",x"1b",x"cd",x"99",x"1e",x"dd",x"71",x"0d",x"dd",x"70",x"0e",
	x"dd",x"36",x"00",x"00",x"2a",x"59",x"5c",x"ed",x"5b",x"53",x"5c",x"37",x"ed",x"52",x"dd",x"75",
	x"0b",x"dd",x"74",x"0c",x"2a",x"4b",x"5c",x"ed",x"52",x"dd",x"75",x"0f",x"dd",x"74",x"10",x"eb",
	x"3a",x"74",x"5c",x"a7",x"ca",x"70",x"09",x"e5",x"01",x"11",x"00",x"dd",x"09",x"dd",x"e5",x"11",
	x"11",x"00",x"af",x"37",x"cd",x"56",x"05",x"dd",x"e1",x"30",x"f2",x"3e",x"fe",x"cd",x"01",x"16",
	x"fd",x"36",x"52",x"03",x"0e",x"80",x"dd",x"7e",x"00",x"dd",x"be",x"ef",x"20",x"02",x"0e",x"f6",
	x"fe",x"04",x"30",x"d9",x"11",x"c0",x"09",x"c5",x"cd",x"0a",x"0c",x"c1",x"dd",x"e5",x"d1",x"21",
	x"f0",x"ff",x"19",x"06",x"0a",x"7e",x"3c",x"20",x"03",x"79",x"80",x"4f",x"13",x"1a",x"be",x"23",
	x"20",x"01",x"0c",x"d7",x"10",x"f6",x"cb",x"79",x"20",x"b3",x"3e",x"0d",x"d7",x"e1",x"dd",x"7e",
	x"00",x"fe",x"03",x"28",x"0c",x"3a",x"74",x"5c",x"3d",x"ca",x"08",x"08",x"fe",x"02",x"ca",x"b6",
	x"08",x"e5",x"dd",x"6e",x"fa",x"dd",x"66",x"fb",x"dd",x"5e",x"0b",x"dd",x"56",x"0c",x"7c",x"b5",
	x"28",x"0d",x"ed",x"52",x"38",x"26",x"28",x"07",x"dd",x"7e",x"00",x"fe",x"03",x"20",x"1d",x"e1",
	x"7c",x"b5",x"20",x"06",x"dd",x"6e",x"0d",x"dd",x"66",x"0e",x"e5",x"dd",x"e1",x"3a",x"74",x"5c",
	x"fe",x"02",x"37",x"20",x"01",x"a7",x"3e",x"ff",x"cd",x"56",x"05",x"d8",x"cf",x"1a",x"dd",x"5e",
	x"0b",x"dd",x"56",x"0c",x"e5",x"7c",x"b5",x"20",x"06",x"13",x"13",x"13",x"eb",x"18",x"0c",x"dd",
	x"6e",x"fa",x"dd",x"66",x"fb",x"eb",x"37",x"ed",x"52",x"38",x"09",x"11",x"05",x"00",x"19",x"44",
	x"4d",x"cd",x"05",x"1f",x"e1",x"dd",x"7e",x"00",x"a7",x"28",x"3e",x"7c",x"b5",x"28",x"13",x"2b",
	x"46",x"2b",x"4e",x"2b",x"03",x"03",x"03",x"dd",x"22",x"5f",x"5c",x"cd",x"e8",x"19",x"dd",x"2a",
	x"5f",x"5c",x"2a",x"59",x"5c",x"2b",x"dd",x"4e",x"0b",x"dd",x"46",x"0c",x"c5",x"03",x"03",x"03",
	x"dd",x"7e",x"fd",x"f5",x"cd",x"55",x"16",x"23",x"f1",x"77",x"d1",x"23",x"73",x"23",x"72",x"23",
	x"e5",x"dd",x"e1",x"37",x"3e",x"ff",x"c3",x"02",x"08",x"eb",x"2a",x"59",x"5c",x"2b",x"dd",x"22",
	x"5f",x"5c",x"dd",x"4e",x"0b",x"dd",x"46",x"0c",x"c5",x"cd",x"e5",x"19",x"c1",x"e5",x"c5",x"cd",
	x"55",x"16",x"dd",x"2a",x"5f",x"5c",x"23",x"dd",x"4e",x"0f",x"dd",x"46",x"10",x"09",x"22",x"4b",
	x"5c",x"dd",x"66",x"0e",x"7c",x"e6",x"c0",x"20",x"0a",x"dd",x"6e",x"0d",x"22",x"42",x"5c",x"fd",
	x"36",x"0a",x"00",x"d1",x"dd",x"e1",x"37",x"3e",x"ff",x"c3",x"02",x"08",x"dd",x"4e",x"0b",x"dd",
	x"46",x"0c",x"c5",x"03",x"f7",x"36",x"80",x"eb",x"d1",x"e5",x"e5",x"dd",x"e1",x"37",x"3e",x"ff",
	x"cd",x"02",x"08",x"e1",x"ed",x"5b",x"53",x"5c",x"7e",x"e6",x"c0",x"20",x"19",x"1a",x"13",x"be",
	x"23",x"20",x"02",x"1a",x"be",x"1b",x"2b",x"30",x"08",x"e5",x"eb",x"cd",x"b8",x"19",x"e1",x"18",
	x"ec",x"cd",x"2c",x"09",x"18",x"e2",x"7e",x"4f",x"fe",x"80",x"c8",x"e5",x"2a",x"4b",x"5c",x"7e",
	x"fe",x"80",x"28",x"25",x"b9",x"28",x"08",x"c5",x"cd",x"b8",x"19",x"c1",x"eb",x"18",x"f0",x"e6",
	x"e0",x"fe",x"a0",x"20",x"12",x"d1",x"d5",x"e5",x"23",x"13",x"1a",x"be",x"20",x"06",x"17",x"30",
	x"f7",x"e1",x"18",x"03",x"e1",x"18",x"e0",x"3e",x"ff",x"d1",x"eb",x"3c",x"37",x"cd",x"2c",x"09",
	x"18",x"c4",x"20",x"10",x"08",x"22",x"5f",x"5c",x"eb",x"cd",x"b8",x"19",x"cd",x"e8",x"19",x"eb",
	x"2a",x"5f",x"5c",x"08",x"08",x"d5",x"cd",x"b8",x"19",x"22",x"5f",x"5c",x"2a",x"53",x"5c",x"e3",
	x"c5",x"08",x"38",x"07",x"2b",x"cd",x"55",x"16",x"23",x"18",x"03",x"cd",x"55",x"16",x"23",x"c1",
	x"d1",x"ed",x"53",x"53",x"5c",x"ed",x"5b",x"5f",x"5c",x"c5",x"d5",x"eb",x"ed",x"b0",x"e1",x"c1",
	x"d5",x"cd",x"e8",x"19",x"d1",x"c9",x"e5",x"3e",x"fd",x"cd",x"01",x"16",x"af",x"11",x"a1",x"09",
	x"cd",x"0a",x"0c",x"fd",x"cb",x"02",x"ee",x"cd",x"d4",x"15",x"dd",x"e5",x"11",x"11",x"00",x"af",
	x"cd",x"c2",x"04",x"dd",x"e1",x"06",x"32",x"76",x"10",x"fd",x"dd",x"5e",x"0b",x"dd",x"56",x"0c",
	x"3e",x"ff",x"dd",x"e1",x"c3",x"c2",x"04",x"80",x"53",x"74",x"61",x"72",x"74",x"20",x"74",x"61",
	x"70",x"65",x"2c",x"20",x"74",x"68",x"65",x"6e",x"20",x"70",x"72",x"65",x"73",x"73",x"20",x"61",
	x"6e",x"79",x"20",x"6b",x"65",x"79",x"ae",x"0d",x"50",x"72",x"6f",x"67",x"72",x"61",x"6d",x"3a",
	x"a0",x"0d",x"4e",x"75",x"6d",x"62",x"65",x"72",x"20",x"61",x"72",x"72",x"61",x"79",x"3a",x"a0",
	x"0d",x"43",x"68",x"61",x"72",x"61",x"63",x"74",x"65",x"72",x"20",x"61",x"72",x"72",x"61",x"79",
	x"3a",x"a0",x"0d",x"42",x"79",x"74",x"65",x"73",x"3a",x"a0",x"cd",x"03",x"0b",x"fe",x"20",x"d2",
	x"d9",x"0a",x"fe",x"06",x"38",x"69",x"fe",x"18",x"30",x"65",x"21",x"0b",x"0a",x"5f",x"16",x"00",
	x"19",x"5e",x"19",x"e5",x"c3",x"03",x"0b",x"4e",x"57",x"10",x"29",x"54",x"53",x"52",x"37",x"50",
	x"4f",x"5f",x"5e",x"5d",x"5c",x"5b",x"5a",x"54",x"53",x"0c",x"3e",x"22",x"b9",x"20",x"11",x"fd",
	x"cb",x"01",x"4e",x"20",x"09",x"04",x"0e",x"02",x"3e",x"18",x"b8",x"20",x"03",x"05",x"0e",x"21",
	x"c3",x"d9",x"0d",x"3a",x"91",x"5c",x"f5",x"fd",x"36",x"57",x"01",x"3e",x"20",x"cd",x"65",x"0b",
	x"f1",x"32",x"91",x"5c",x"c9",x"fd",x"cb",x"01",x"4e",x"c2",x"cd",x"0e",x"0e",x"21",x"cd",x"55",
	x"0c",x"05",x"c3",x"d9",x"0d",x"cd",x"03",x"0b",x"79",x"3d",x"3d",x"e6",x"10",x"18",x"5a",x"3e",
	x"3f",x"18",x"6c",x"11",x"87",x"0a",x"32",x"0f",x"5c",x"18",x"0b",x"11",x"6d",x"0a",x"18",x"03",
	x"11",x"87",x"0a",x"32",x"0e",x"5c",x"2a",x"51",x"5c",x"73",x"23",x"72",x"c9",x"11",x"f4",x"09",
	x"cd",x"80",x"0a",x"2a",x"0e",x"5c",x"57",x"7d",x"fe",x"16",x"da",x"11",x"22",x"20",x"29",x"44",
	x"4a",x"3e",x"1f",x"91",x"38",x"0c",x"c6",x"02",x"4f",x"fd",x"cb",x"01",x"4e",x"20",x"16",x"3e",
	x"16",x"90",x"da",x"9f",x"1e",x"3c",x"47",x"04",x"fd",x"cb",x"02",x"46",x"c2",x"55",x"0c",x"fd",
	x"be",x"31",x"da",x"86",x"0c",x"c3",x"d9",x"0d",x"7c",x"cd",x"03",x"0b",x"81",x"3d",x"e6",x"1f",
	x"c8",x"57",x"fd",x"cb",x"01",x"c6",x"3e",x"20",x"cd",x"3b",x"0c",x"15",x"20",x"f8",x"c9",x"cd",
	x"24",x"0b",x"fd",x"cb",x"01",x"4e",x"20",x"1a",x"fd",x"cb",x"02",x"46",x"20",x"08",x"ed",x"43",
	x"88",x"5c",x"22",x"84",x"5c",x"c9",x"ed",x"43",x"8a",x"5c",x"ed",x"43",x"82",x"5c",x"22",x"86",
	x"5c",x"c9",x"fd",x"71",x"45",x"22",x"80",x"5c",x"c9",x"fd",x"cb",x"01",x"4e",x"20",x"14",x"ed",
	x"4b",x"88",x"5c",x"2a",x"84",x"5c",x"fd",x"cb",x"02",x"46",x"c8",x"ed",x"4b",x"8a",x"5c",x"2a",
	x"86",x"5c",x"c9",x"fd",x"4e",x"45",x"2a",x"80",x"5c",x"c9",x"fe",x"80",x"38",x"3d",x"fe",x"90",
	x"30",x"26",x"47",x"cd",x"38",x"0b",x"cd",x"03",x"0b",x"11",x"92",x"5c",x"18",x"47",x"21",x"92",
	x"5c",x"cd",x"3e",x"0b",x"cb",x"18",x"9f",x"e6",x"0f",x"4f",x"cb",x"18",x"9f",x"e6",x"f0",x"b1",
	x"0e",x"04",x"77",x"23",x"0d",x"20",x"fb",x"c9",x"d6",x"a5",x"30",x"09",x"c6",x"15",x"c5",x"ed",
	x"4b",x"7b",x"5c",x"18",x"0b",x"cd",x"10",x"0c",x"c3",x"03",x"0b",x"c5",x"ed",x"4b",x"36",x"5c",
	x"eb",x"21",x"3b",x"5c",x"cb",x"86",x"fe",x"20",x"20",x"02",x"cb",x"c6",x"26",x"00",x"6f",x"29",
	x"29",x"29",x"09",x"c1",x"eb",x"79",x"3d",x"3e",x"21",x"20",x"0e",x"05",x"4f",x"fd",x"cb",x"01",
	x"4e",x"28",x"06",x"d5",x"cd",x"cd",x"0e",x"d1",x"79",x"b9",x"d5",x"cc",x"55",x"0c",x"d1",x"c5",
	x"e5",x"3a",x"91",x"5c",x"06",x"ff",x"1f",x"38",x"01",x"04",x"1f",x"1f",x"9f",x"4f",x"3e",x"08",
	x"a7",x"fd",x"cb",x"01",x"4e",x"28",x"05",x"fd",x"cb",x"30",x"ce",x"37",x"eb",x"08",x"1a",x"a0",
	x"ae",x"a9",x"12",x"08",x"38",x"13",x"14",x"23",x"3d",x"20",x"f2",x"eb",x"25",x"fd",x"cb",x"01",
	x"4e",x"cc",x"db",x"0b",x"e1",x"c1",x"0d",x"23",x"c9",x"08",x"3e",x"20",x"83",x"5f",x"08",x"18",
	x"e6",x"7c",x"0f",x"0f",x"0f",x"e6",x"03",x"f6",x"58",x"67",x"ed",x"5b",x"8f",x"5c",x"7e",x"ab",
	x"a2",x"ab",x"fd",x"cb",x"57",x"76",x"28",x"08",x"e6",x"c7",x"cb",x"57",x"20",x"02",x"ee",x"38",
	x"fd",x"cb",x"57",x"66",x"28",x"08",x"e6",x"f8",x"cb",x"6f",x"20",x"02",x"ee",x"07",x"77",x"c9",
	x"e5",x"26",x"00",x"e3",x"18",x"04",x"11",x"95",x"00",x"f5",x"cd",x"41",x"0c",x"38",x"09",x"3e",
	x"20",x"fd",x"cb",x"01",x"46",x"cc",x"3b",x"0c",x"1a",x"e6",x"7f",x"cd",x"3b",x"0c",x"1a",x"13",
	x"87",x"30",x"f5",x"d1",x"fe",x"48",x"28",x"03",x"fe",x"82",x"d8",x"7a",x"fe",x"03",x"d8",x"3e",
	x"20",x"d5",x"d9",x"d7",x"d9",x"d1",x"c9",x"f5",x"eb",x"3c",x"cb",x"7e",x"23",x"28",x"fb",x"3d",
	x"20",x"f8",x"eb",x"f1",x"fe",x"20",x"d8",x"1a",x"d6",x"41",x"c9",x"fd",x"cb",x"01",x"4e",x"c0",
	x"11",x"d9",x"0d",x"d5",x"78",x"fd",x"cb",x"02",x"46",x"c2",x"02",x"0d",x"fd",x"be",x"31",x"38",
	x"1b",x"c0",x"fd",x"cb",x"02",x"66",x"28",x"16",x"fd",x"5e",x"2d",x"1d",x"28",x"5a",x"3e",x"00",
	x"cd",x"01",x"16",x"ed",x"7b",x"3f",x"5c",x"fd",x"cb",x"02",x"a6",x"c9",x"cf",x"04",x"fd",x"35",
	x"52",x"20",x"45",x"3e",x"18",x"90",x"32",x"8c",x"5c",x"2a",x"8f",x"5c",x"e5",x"3a",x"91",x"5c",
	x"f5",x"3e",x"fd",x"cd",x"01",x"16",x"af",x"11",x"f8",x"0c",x"cd",x"0a",x"0c",x"fd",x"cb",x"02",
	x"ee",x"21",x"3b",x"5c",x"cb",x"de",x"cb",x"ae",x"d9",x"cd",x"d4",x"15",x"d9",x"fe",x"20",x"28",
	x"45",x"fe",x"e2",x"28",x"41",x"f6",x"20",x"fe",x"6e",x"28",x"3b",x"3e",x"fe",x"cd",x"01",x"16",
	x"f1",x"32",x"91",x"5c",x"e1",x"22",x"8f",x"5c",x"cd",x"fe",x"0d",x"fd",x"46",x"31",x"04",x"0e",
	x"21",x"c5",x"cd",x"9b",x"0e",x"7c",x"0f",x"0f",x"0f",x"e6",x"03",x"f6",x"58",x"67",x"11",x"e0",
	x"5a",x"1a",x"4e",x"06",x"20",x"eb",x"12",x"71",x"13",x"23",x"10",x"fa",x"c1",x"c9",x"80",x"73",
	x"63",x"72",x"6f",x"6c",x"6c",x"bf",x"cf",x"0c",x"fe",x"02",x"38",x"80",x"fd",x"86",x"31",x"d6",
	x"19",x"d0",x"ed",x"44",x"c5",x"47",x"2a",x"8f",x"5c",x"e5",x"2a",x"91",x"5c",x"e5",x"cd",x"4d",
	x"0d",x"78",x"f5",x"21",x"6b",x"5c",x"46",x"78",x"3c",x"77",x"21",x"89",x"5c",x"be",x"38",x"03",
	x"34",x"06",x"18",x"cd",x"00",x"0e",x"f1",x"3d",x"20",x"e8",x"e1",x"fd",x"75",x"57",x"e1",x"22",
	x"8f",x"5c",x"ed",x"4b",x"88",x"5c",x"fd",x"cb",x"02",x"86",x"cd",x"d9",x"0d",x"fd",x"cb",x"02",
	x"c6",x"c1",x"c9",x"af",x"2a",x"8d",x"5c",x"fd",x"cb",x"02",x"46",x"28",x"04",x"67",x"fd",x"6e",
	x"0e",x"22",x"8f",x"5c",x"21",x"91",x"5c",x"20",x"02",x"7e",x"0f",x"ae",x"e6",x"55",x"ae",x"77",
	x"c9",x"cd",x"af",x"0d",x"21",x"3c",x"5c",x"cb",x"ae",x"cb",x"c6",x"cd",x"4d",x"0d",x"fd",x"46",
	x"31",x"cd",x"44",x"0e",x"21",x"c0",x"5a",x"3a",x"8d",x"5c",x"05",x"18",x"07",x"0e",x"20",x"2b",
	x"77",x"0d",x"20",x"fb",x"10",x"f7",x"fd",x"36",x"31",x"02",x"3e",x"fd",x"cd",x"01",x"16",x"2a",
	x"51",x"5c",x"11",x"f4",x"09",x"a7",x"73",x"23",x"72",x"23",x"11",x"a8",x"10",x"3f",x"38",x"f6",
	x"01",x"21",x"17",x"18",x"2a",x"21",x"00",x"00",x"22",x"7d",x"5c",x"fd",x"cb",x"30",x"86",x"cd",
	x"94",x"0d",x"3e",x"fe",x"cd",x"01",x"16",x"cd",x"4d",x"0d",x"06",x"18",x"cd",x"44",x"0e",x"2a",
	x"51",x"5c",x"11",x"f4",x"09",x"73",x"23",x"72",x"fd",x"36",x"52",x"01",x"01",x"21",x"18",x"21",
	x"00",x"5b",x"fd",x"cb",x"01",x"4e",x"20",x"12",x"78",x"fd",x"cb",x"02",x"46",x"28",x"05",x"fd",
	x"86",x"31",x"d6",x"18",x"c5",x"47",x"cd",x"9b",x"0e",x"c1",x"3e",x"21",x"91",x"5f",x"16",x"00",
	x"19",x"c3",x"dc",x"0a",x"06",x"17",x"cd",x"9b",x"0e",x"0e",x"08",x"c5",x"e5",x"78",x"e6",x"07",
	x"78",x"20",x"0c",x"eb",x"21",x"e0",x"f8",x"19",x"eb",x"01",x"20",x"00",x"3d",x"ed",x"b0",x"eb",
	x"21",x"e0",x"ff",x"19",x"eb",x"47",x"e6",x"07",x"0f",x"0f",x"0f",x"4f",x"78",x"06",x"00",x"ed",
	x"b0",x"06",x"07",x"09",x"e6",x"f8",x"20",x"db",x"e1",x"24",x"c1",x"0d",x"20",x"cd",x"cd",x"88",
	x"0e",x"21",x"e0",x"ff",x"19",x"eb",x"ed",x"b0",x"06",x"01",x"c5",x"cd",x"9b",x"0e",x"0e",x"08",
	x"c5",x"e5",x"78",x"e6",x"07",x"0f",x"0f",x"0f",x"4f",x"78",x"06",x"00",x"0d",x"54",x"5d",x"36",
	x"00",x"13",x"ed",x"b0",x"11",x"01",x"07",x"19",x"3d",x"e6",x"f8",x"47",x"20",x"e5",x"e1",x"24",
	x"c1",x"0d",x"20",x"dc",x"cd",x"88",x"0e",x"62",x"6b",x"13",x"3a",x"8d",x"5c",x"fd",x"cb",x"02",
	x"46",x"28",x"03",x"3a",x"48",x"5c",x"77",x"0b",x"ed",x"b0",x"c1",x"0e",x"21",x"c9",x"7c",x"0f",
	x"0f",x"0f",x"3d",x"f6",x"50",x"67",x"eb",x"61",x"68",x"29",x"29",x"29",x"29",x"29",x"44",x"4d",
	x"c9",x"3e",x"18",x"90",x"57",x"0f",x"0f",x"0f",x"e6",x"e0",x"6f",x"7a",x"e6",x"18",x"f6",x"40",
	x"67",x"c9",x"f3",x"06",x"b0",x"21",x"00",x"40",x"e5",x"c5",x"cd",x"f4",x"0e",x"c1",x"e1",x"24",
	x"7c",x"e6",x"07",x"20",x"0a",x"7d",x"c6",x"20",x"6f",x"3f",x"9f",x"e6",x"f8",x"84",x"67",x"10",
	x"e7",x"18",x"0d",x"f3",x"21",x"00",x"5b",x"06",x"08",x"c5",x"cd",x"f4",x"0e",x"c1",x"10",x"f9",
	x"3e",x"04",x"d3",x"fb",x"fb",x"21",x"00",x"5b",x"fd",x"75",x"46",x"af",x"47",x"77",x"23",x"10",
	x"fc",x"fd",x"cb",x"30",x"8e",x"0e",x"21",x"c3",x"d9",x"0d",x"78",x"fe",x"03",x"9f",x"e6",x"02",
	x"d3",x"fb",x"57",x"cd",x"54",x"1f",x"38",x"0a",x"3e",x"04",x"d3",x"fb",x"fb",x"cd",x"df",x"0e",
	x"cf",x"0c",x"db",x"fb",x"87",x"f8",x"30",x"eb",x"0e",x"20",x"5e",x"23",x"06",x"08",x"cb",x"12",
	x"cb",x"13",x"cb",x"1a",x"db",x"fb",x"1f",x"30",x"fb",x"7a",x"d3",x"fb",x"10",x"f0",x"0d",x"20",
	x"e9",x"c9",x"2a",x"3d",x"5c",x"e5",x"21",x"7f",x"10",x"e5",x"ed",x"73",x"3d",x"5c",x"cd",x"d4",
	x"15",x"f5",x"16",x"00",x"fd",x"5e",x"ff",x"21",x"c8",x"00",x"cd",x"b5",x"03",x"f1",x"21",x"38",
	x"0f",x"e5",x"fe",x"18",x"30",x"31",x"fe",x"07",x"38",x"2d",x"fe",x"10",x"38",x"3a",x"01",x"02",
	x"00",x"57",x"fe",x"16",x"38",x"0c",x"03",x"fd",x"cb",x"37",x"7e",x"ca",x"1e",x"10",x"cd",x"d4",
	x"15",x"5f",x"cd",x"d4",x"15",x"d5",x"2a",x"5b",x"5c",x"fd",x"cb",x"07",x"86",x"cd",x"55",x"16",
	x"c1",x"23",x"70",x"23",x"71",x"18",x"0a",x"fd",x"cb",x"07",x"86",x"2a",x"5b",x"5c",x"cd",x"52",
	x"16",x"12",x"13",x"ed",x"53",x"5b",x"5c",x"c9",x"5f",x"16",x"00",x"21",x"99",x"0f",x"19",x"5e",
	x"19",x"e5",x"2a",x"5b",x"5c",x"c9",x"09",x"66",x"6a",x"50",x"b5",x"70",x"7e",x"cf",x"d4",x"2a",
	x"49",x"5c",x"fd",x"cb",x"37",x"6e",x"c2",x"97",x"10",x"cd",x"6e",x"19",x"cd",x"95",x"16",x"7a",
	x"b3",x"ca",x"97",x"10",x"e5",x"23",x"4e",x"23",x"46",x"21",x"0a",x"00",x"09",x"44",x"4d",x"cd",
	x"05",x"1f",x"cd",x"97",x"10",x"2a",x"51",x"5c",x"e3",x"e5",x"3e",x"ff",x"cd",x"01",x"16",x"e1",
	x"2b",x"fd",x"35",x"0f",x"cd",x"55",x"18",x"fd",x"34",x"0f",x"2a",x"59",x"5c",x"23",x"23",x"23",
	x"23",x"22",x"5b",x"5c",x"e1",x"cd",x"15",x"16",x"c9",x"fd",x"cb",x"37",x"6e",x"20",x"08",x"21",
	x"49",x"5c",x"cd",x"0f",x"19",x"18",x"6d",x"fd",x"36",x"00",x"10",x"18",x"1d",x"cd",x"31",x"10",
	x"18",x"05",x"7e",x"fe",x"0d",x"c8",x"23",x"22",x"5b",x"5c",x"c9",x"cd",x"31",x"10",x"01",x"01",
	x"00",x"c3",x"e8",x"19",x"cd",x"d4",x"15",x"cd",x"d4",x"15",x"e1",x"e1",x"e1",x"22",x"3d",x"5c",
	x"fd",x"cb",x"00",x"7e",x"c0",x"f9",x"c9",x"37",x"cd",x"95",x"11",x"ed",x"52",x"19",x"23",x"c1",
	x"d8",x"c5",x"44",x"4d",x"62",x"6b",x"23",x"1a",x"e6",x"f0",x"fe",x"10",x"20",x"09",x"23",x"1a",
	x"d6",x"17",x"ce",x"00",x"20",x"01",x"23",x"a7",x"ed",x"42",x"09",x"eb",x"38",x"e6",x"c9",x"fd",
	x"cb",x"37",x"6e",x"c0",x"2a",x"49",x"5c",x"cd",x"6e",x"19",x"eb",x"cd",x"95",x"16",x"21",x"4a",
	x"5c",x"cd",x"1c",x"19",x"cd",x"95",x"17",x"3e",x"00",x"c3",x"01",x"16",x"fd",x"cb",x"37",x"7e",
	x"28",x"a8",x"c3",x"81",x"0f",x"fd",x"cb",x"30",x"66",x"28",x"a1",x"fd",x"36",x"00",x"ff",x"16",
	x"00",x"fd",x"5e",x"fe",x"21",x"90",x"1a",x"cd",x"b5",x"03",x"c3",x"30",x"0f",x"e5",x"cd",x"90",
	x"11",x"2b",x"cd",x"e5",x"19",x"22",x"5b",x"5c",x"fd",x"36",x"07",x"00",x"e1",x"c9",x"fd",x"cb",
	x"02",x"5e",x"c4",x"1d",x"11",x"a7",x"fd",x"cb",x"01",x"6e",x"c8",x"3a",x"08",x"5c",x"fd",x"cb",
	x"01",x"ae",x"f5",x"fd",x"cb",x"02",x"6e",x"c4",x"6e",x"0d",x"f1",x"fe",x"20",x"30",x"52",x"fe",
	x"10",x"30",x"2d",x"fe",x"06",x"30",x"0a",x"47",x"e6",x"01",x"4f",x"78",x"1f",x"c6",x"12",x"18",
	x"2a",x"20",x"09",x"21",x"6a",x"5c",x"3e",x"08",x"ae",x"77",x"18",x"0e",x"fe",x"0e",x"d8",x"d6",
	x"0d",x"21",x"41",x"5c",x"be",x"77",x"20",x"02",x"36",x"00",x"fd",x"cb",x"02",x"de",x"bf",x"c9",
	x"47",x"e6",x"07",x"4f",x"3e",x"10",x"cb",x"58",x"20",x"01",x"3c",x"fd",x"71",x"d3",x"11",x"0d",
	x"11",x"18",x"06",x"3a",x"0d",x"5c",x"11",x"a8",x"10",x"2a",x"4f",x"5c",x"23",x"23",x"73",x"23",
	x"72",x"37",x"c9",x"cd",x"4d",x"0d",x"fd",x"cb",x"02",x"9e",x"fd",x"cb",x"02",x"ae",x"2a",x"8a",
	x"5c",x"e5",x"2a",x"3d",x"5c",x"e5",x"21",x"67",x"11",x"e5",x"ed",x"73",x"3d",x"5c",x"2a",x"82",
	x"5c",x"e5",x"37",x"cd",x"95",x"11",x"eb",x"cd",x"7d",x"18",x"eb",x"cd",x"e1",x"18",x"2a",x"8a",
	x"5c",x"e3",x"eb",x"cd",x"4d",x"0d",x"3a",x"8b",x"5c",x"92",x"38",x"26",x"20",x"06",x"7b",x"fd",
	x"96",x"50",x"30",x"1e",x"3e",x"20",x"d5",x"cd",x"f4",x"09",x"d1",x"18",x"e9",x"16",x"00",x"fd",
	x"5e",x"fe",x"21",x"90",x"1a",x"cd",x"b5",x"03",x"fd",x"36",x"00",x"ff",x"ed",x"5b",x"8a",x"5c",
	x"18",x"02",x"d1",x"e1",x"e1",x"22",x"3d",x"5c",x"c1",x"d5",x"cd",x"d9",x"0d",x"e1",x"22",x"82",
	x"5c",x"fd",x"36",x"26",x"00",x"c9",x"2a",x"61",x"5c",x"2b",x"a7",x"ed",x"5b",x"59",x"5c",x"fd",
	x"cb",x"37",x"6e",x"c8",x"ed",x"5b",x"61",x"5c",x"d8",x"2a",x"63",x"5c",x"c9",x"7e",x"fe",x"0e",
	x"01",x"06",x"00",x"cc",x"e8",x"19",x"7e",x"23",x"fe",x"0d",x"20",x"f1",x"c9",x"f3",x"3e",x"ff",
	x"ed",x"5b",x"b2",x"5c",x"d9",x"ed",x"4b",x"b4",x"5c",x"ed",x"5b",x"38",x"5c",x"2a",x"7b",x"5c",
	x"d9",x"47",x"3e",x"07",x"d3",x"fe",x"3e",x"3f",x"ed",x"47",x"00",x"00",x"00",x"00",x"00",x"00",
	x"62",x"6b",x"36",x"02",x"2b",x"bc",x"20",x"fa",x"a7",x"ed",x"52",x"19",x"23",x"30",x"06",x"35",
	x"28",x"03",x"35",x"28",x"f3",x"2b",x"d9",x"ed",x"43",x"b4",x"5c",x"ed",x"53",x"38",x"5c",x"22",
	x"7b",x"5c",x"d9",x"04",x"28",x"19",x"22",x"b4",x"5c",x"11",x"af",x"3e",x"01",x"a8",x"00",x"eb",
	x"ed",x"b8",x"eb",x"23",x"22",x"7b",x"5c",x"2b",x"01",x"40",x"00",x"ed",x"43",x"38",x"5c",x"22",
	x"b2",x"5c",x"21",x"00",x"3c",x"22",x"36",x"5c",x"2a",x"b2",x"5c",x"36",x"3e",x"2b",x"f9",x"2b",
	x"2b",x"22",x"3d",x"5c",x"ed",x"56",x"fd",x"21",x"3a",x"5c",x"fb",x"21",x"b6",x"5c",x"22",x"4f",
	x"5c",x"11",x"af",x"15",x"01",x"15",x"00",x"eb",x"ed",x"b0",x"eb",x"2b",x"22",x"57",x"5c",x"23",
	x"22",x"53",x"5c",x"22",x"4b",x"5c",x"36",x"80",x"23",x"22",x"59",x"5c",x"36",x"0d",x"23",x"36",
	x"80",x"23",x"22",x"61",x"5c",x"22",x"63",x"5c",x"22",x"65",x"5c",x"3e",x"38",x"32",x"8d",x"5c",
	x"32",x"8f",x"5c",x"32",x"48",x"5c",x"21",x"23",x"05",x"22",x"09",x"5c",x"fd",x"35",x"c6",x"fd",
	x"35",x"ca",x"21",x"c6",x"15",x"11",x"10",x"5c",x"01",x"0e",x"00",x"ed",x"b0",x"fd",x"cb",x"01",
	x"ce",x"cd",x"df",x"0e",x"fd",x"36",x"31",x"02",x"cd",x"6b",x"0d",x"af",x"11",x"38",x"15",x"cd",
	x"0a",x"0c",x"fd",x"cb",x"02",x"ee",x"18",x"07",x"fd",x"36",x"31",x"02",x"cd",x"95",x"17",x"cd",
	x"b0",x"16",x"3e",x"00",x"cd",x"01",x"16",x"cd",x"2c",x"0f",x"cd",x"17",x"1b",x"fd",x"cb",x"00",
	x"7e",x"20",x"12",x"fd",x"cb",x"30",x"66",x"28",x"40",x"2a",x"59",x"5c",x"cd",x"a7",x"11",x"fd",
	x"36",x"00",x"ff",x"18",x"dd",x"2a",x"59",x"5c",x"22",x"5d",x"5c",x"cd",x"fb",x"19",x"78",x"b1",
	x"c2",x"5d",x"15",x"df",x"fe",x"0d",x"28",x"c0",x"fd",x"cb",x"30",x"46",x"c4",x"af",x"0d",x"cd",
	x"6e",x"0d",x"3e",x"19",x"fd",x"96",x"4f",x"32",x"8c",x"5c",x"fd",x"cb",x"01",x"fe",x"fd",x"36",
	x"00",x"ff",x"fd",x"36",x"0a",x"01",x"cd",x"8a",x"1b",x"76",x"fd",x"cb",x"01",x"ae",x"fd",x"cb",
	x"30",x"4e",x"c4",x"cd",x"0e",x"3a",x"3a",x"5c",x"3c",x"f5",x"21",x"00",x"00",x"fd",x"74",x"37",
	x"fd",x"74",x"26",x"22",x"0b",x"5c",x"21",x"01",x"00",x"22",x"16",x"5c",x"cd",x"b0",x"16",x"fd",
	x"cb",x"37",x"ae",x"cd",x"6e",x"0d",x"fd",x"cb",x"02",x"ee",x"f1",x"47",x"fe",x"0a",x"38",x"02",
	x"c6",x"07",x"cd",x"ef",x"15",x"3e",x"20",x"d7",x"78",x"11",x"91",x"13",x"cd",x"0a",x"0c",x"af",
	x"11",x"36",x"15",x"cd",x"0a",x"0c",x"ed",x"4b",x"45",x"5c",x"cd",x"1b",x"1a",x"3e",x"3a",x"d7",
	x"fd",x"4e",x"0d",x"06",x"00",x"cd",x"1b",x"1a",x"cd",x"97",x"10",x"3a",x"3a",x"5c",x"3c",x"28",
	x"1b",x"fe",x"09",x"28",x"04",x"fe",x"15",x"20",x"03",x"fd",x"34",x"0d",x"01",x"03",x"00",x"11",
	x"70",x"5c",x"21",x"44",x"5c",x"cb",x"7e",x"28",x"01",x"09",x"ed",x"b8",x"fd",x"36",x"0a",x"ff",
	x"fd",x"cb",x"01",x"9e",x"c3",x"ac",x"12",x"80",x"4f",x"cb",x"4e",x"45",x"58",x"54",x"20",x"77",
	x"69",x"74",x"68",x"6f",x"75",x"74",x"20",x"46",x"4f",x"d2",x"56",x"61",x"72",x"69",x"61",x"62",
	x"6c",x"65",x"20",x"6e",x"6f",x"74",x"20",x"66",x"6f",x"75",x"6e",x"e4",x"53",x"75",x"62",x"73",
	x"63",x"72",x"69",x"70",x"74",x"20",x"77",x"72",x"6f",x"6e",x"e7",x"4f",x"75",x"74",x"20",x"6f",
	x"66",x"20",x"6d",x"65",x"6d",x"6f",x"72",x"f9",x"4f",x"75",x"74",x"20",x"6f",x"66",x"20",x"73",
	x"63",x"72",x"65",x"65",x"ee",x"4e",x"75",x"6d",x"62",x"65",x"72",x"20",x"74",x"6f",x"6f",x"20",
	x"62",x"69",x"e7",x"52",x"45",x"54",x"55",x"52",x"4e",x"20",x"77",x"69",x"74",x"68",x"6f",x"75",
	x"74",x"20",x"47",x"4f",x"53",x"55",x"c2",x"45",x"6e",x"64",x"20",x"6f",x"66",x"20",x"66",x"69",
	x"6c",x"e5",x"53",x"54",x"4f",x"50",x"20",x"73",x"74",x"61",x"74",x"65",x"6d",x"65",x"6e",x"f4",
	x"49",x"6e",x"76",x"61",x"6c",x"69",x"64",x"20",x"61",x"72",x"67",x"75",x"6d",x"65",x"6e",x"f4",
	x"49",x"6e",x"74",x"65",x"67",x"65",x"72",x"20",x"6f",x"75",x"74",x"20",x"6f",x"66",x"20",x"72",
	x"61",x"6e",x"67",x"e5",x"4e",x"6f",x"6e",x"73",x"65",x"6e",x"73",x"65",x"20",x"69",x"6e",x"20",
	x"42",x"41",x"53",x"49",x"c3",x"42",x"52",x"45",x"41",x"4b",x"20",x"2d",x"20",x"43",x"4f",x"4e",
	x"54",x"20",x"72",x"65",x"70",x"65",x"61",x"74",x"f3",x"4f",x"75",x"74",x"20",x"6f",x"66",x"20",
	x"44",x"41",x"54",x"c1",x"49",x"6e",x"76",x"61",x"6c",x"69",x"64",x"20",x"66",x"69",x"6c",x"65",
	x"20",x"6e",x"61",x"6d",x"e5",x"4e",x"6f",x"20",x"72",x"6f",x"6f",x"6d",x"20",x"66",x"6f",x"72",
	x"20",x"6c",x"69",x"6e",x"e5",x"53",x"54",x"4f",x"50",x"20",x"69",x"6e",x"20",x"49",x"4e",x"50",
	x"55",x"d4",x"46",x"4f",x"52",x"20",x"77",x"69",x"74",x"68",x"6f",x"75",x"74",x"20",x"4e",x"45",
	x"58",x"d4",x"49",x"6e",x"76",x"61",x"6c",x"69",x"64",x"20",x"49",x"2f",x"4f",x"20",x"64",x"65",
	x"76",x"69",x"63",x"e5",x"49",x"6e",x"76",x"61",x"6c",x"69",x"64",x"20",x"63",x"6f",x"6c",x"6f",
	x"75",x"f2",x"42",x"52",x"45",x"41",x"4b",x"20",x"69",x"6e",x"74",x"6f",x"20",x"70",x"72",x"6f",
	x"67",x"72",x"61",x"ed",x"52",x"41",x"4d",x"54",x"4f",x"50",x"20",x"6e",x"6f",x"20",x"67",x"6f",
	x"6f",x"e4",x"53",x"74",x"61",x"74",x"65",x"6d",x"65",x"6e",x"74",x"20",x"6c",x"6f",x"73",x"f4",
	x"49",x"6e",x"76",x"61",x"6c",x"69",x"64",x"20",x"73",x"74",x"72",x"65",x"61",x"ed",x"46",x"4e",
	x"20",x"77",x"69",x"74",x"68",x"6f",x"75",x"74",x"20",x"44",x"45",x"c6",x"50",x"61",x"72",x"61",
	x"6d",x"65",x"74",x"65",x"72",x"20",x"65",x"72",x"72",x"6f",x"f2",x"54",x"61",x"70",x"65",x"20",
	x"6c",x"6f",x"61",x"64",x"69",x"6e",x"67",x"20",x"65",x"72",x"72",x"6f",x"f2",x"2c",x"a0",x"7f",
	x"20",x"31",x"39",x"38",x"32",x"20",x"53",x"69",x"6e",x"63",x"6c",x"61",x"69",x"72",x"20",x"52",
	x"65",x"73",x"65",x"61",x"72",x"63",x"68",x"20",x"4c",x"74",x"e4",x"3e",x"10",x"01",x"00",x"00",
	x"c3",x"13",x"13",x"ed",x"43",x"49",x"5c",x"2a",x"5d",x"5c",x"eb",x"21",x"55",x"15",x"e5",x"2a",
	x"61",x"5c",x"37",x"ed",x"52",x"e5",x"60",x"69",x"cd",x"6e",x"19",x"20",x"06",x"cd",x"b8",x"19",
	x"cd",x"e8",x"19",x"c1",x"79",x"3d",x"b0",x"28",x"28",x"c5",x"03",x"03",x"03",x"03",x"2b",x"ed",
	x"5b",x"53",x"5c",x"d5",x"cd",x"55",x"16",x"e1",x"22",x"53",x"5c",x"c1",x"c5",x"13",x"2a",x"61",
	x"5c",x"2b",x"2b",x"ed",x"b8",x"2a",x"49",x"5c",x"eb",x"c1",x"70",x"2b",x"71",x"2b",x"73",x"2b",
	x"72",x"f1",x"c3",x"a2",x"12",x"f4",x"09",x"a8",x"10",x"4b",x"f4",x"09",x"c4",x"15",x"53",x"81",
	x"0f",x"c4",x"15",x"52",x"f4",x"09",x"c4",x"15",x"50",x"80",x"cf",x"12",x"01",x"00",x"06",x"00",
	x"0b",x"00",x"01",x"00",x"01",x"00",x"06",x"00",x"10",x"00",x"fd",x"cb",x"02",x"6e",x"20",x"04",
	x"fd",x"cb",x"02",x"de",x"cd",x"e6",x"15",x"d8",x"28",x"fa",x"cf",x"07",x"d9",x"e5",x"2a",x"51",
	x"5c",x"23",x"23",x"18",x"08",x"1e",x"30",x"83",x"d9",x"e5",x"2a",x"51",x"5c",x"5e",x"23",x"56",
	x"eb",x"cd",x"2c",x"16",x"e1",x"d9",x"c9",x"87",x"c6",x"16",x"6f",x"26",x"5c",x"5e",x"23",x"56",
	x"7a",x"b3",x"20",x"02",x"cf",x"17",x"1b",x"2a",x"4f",x"5c",x"19",x"22",x"51",x"5c",x"fd",x"cb",
	x"30",x"a6",x"23",x"23",x"23",x"23",x"4e",x"21",x"2d",x"16",x"cd",x"dc",x"16",x"d0",x"16",x"00",
	x"5e",x"19",x"e9",x"4b",x"06",x"53",x"12",x"50",x"1b",x"00",x"fd",x"cb",x"02",x"c6",x"fd",x"cb",
	x"01",x"ae",x"fd",x"cb",x"30",x"e6",x"18",x"04",x"fd",x"cb",x"02",x"86",x"fd",x"cb",x"01",x"8e",
	x"c3",x"4d",x"0d",x"fd",x"cb",x"01",x"ce",x"c9",x"01",x"01",x"00",x"e5",x"cd",x"05",x"1f",x"e1",
	x"cd",x"64",x"16",x"2a",x"65",x"5c",x"eb",x"ed",x"b8",x"c9",x"f5",x"e5",x"21",x"4b",x"5c",x"3e",
	x"0e",x"5e",x"23",x"56",x"e3",x"a7",x"ed",x"52",x"19",x"e3",x"30",x"09",x"d5",x"eb",x"09",x"eb",
	x"72",x"2b",x"73",x"23",x"d1",x"23",x"3d",x"20",x"e8",x"eb",x"d1",x"f1",x"a7",x"ed",x"52",x"44",
	x"4d",x"03",x"19",x"eb",x"c9",x"00",x"00",x"eb",x"11",x"8f",x"16",x"7e",x"e6",x"c0",x"20",x"f7",
	x"56",x"23",x"5e",x"c9",x"2a",x"63",x"5c",x"2b",x"cd",x"55",x"16",x"23",x"23",x"c1",x"ed",x"43",
	x"61",x"5c",x"c1",x"eb",x"23",x"c9",x"2a",x"59",x"5c",x"36",x"0d",x"22",x"5b",x"5c",x"23",x"36",
	x"80",x"23",x"22",x"61",x"5c",x"2a",x"61",x"5c",x"22",x"63",x"5c",x"2a",x"63",x"5c",x"22",x"65",
	x"5c",x"e5",x"21",x"92",x"5c",x"22",x"68",x"5c",x"e1",x"c9",x"ed",x"5b",x"59",x"5c",x"c3",x"e5",
	x"19",x"23",x"7e",x"a7",x"c8",x"b9",x"23",x"20",x"f8",x"37",x"c9",x"cd",x"1e",x"17",x"cd",x"01",
	x"17",x"01",x"00",x"00",x"11",x"e2",x"a3",x"eb",x"19",x"38",x"07",x"01",x"d4",x"15",x"09",x"4e",
	x"23",x"46",x"eb",x"71",x"23",x"70",x"c9",x"e5",x"2a",x"4f",x"5c",x"09",x"23",x"23",x"23",x"4e",
	x"eb",x"21",x"16",x"17",x"cd",x"dc",x"16",x"4e",x"06",x"00",x"09",x"e9",x"4b",x"05",x"53",x"03",
	x"50",x"01",x"e1",x"c9",x"cd",x"94",x"1e",x"fe",x"10",x"38",x"02",x"cf",x"17",x"c6",x"03",x"07",
	x"21",x"10",x"5c",x"4f",x"06",x"00",x"09",x"4e",x"23",x"46",x"2b",x"c9",x"ef",x"01",x"38",x"cd",
	x"1e",x"17",x"78",x"b1",x"28",x"16",x"eb",x"2a",x"4f",x"5c",x"09",x"23",x"23",x"23",x"7e",x"eb",
	x"fe",x"4b",x"28",x"08",x"fe",x"53",x"28",x"04",x"fe",x"50",x"20",x"cf",x"cd",x"5d",x"17",x"73",
	x"23",x"72",x"c9",x"e5",x"cd",x"f1",x"2b",x"78",x"b1",x"20",x"02",x"cf",x"0e",x"c5",x"1a",x"e6",
	x"df",x"4f",x"21",x"7a",x"17",x"cd",x"dc",x"16",x"30",x"f1",x"4e",x"06",x"00",x"09",x"c1",x"e9",
	x"4b",x"06",x"53",x"08",x"50",x"0a",x"00",x"1e",x"01",x"18",x"06",x"1e",x"06",x"18",x"02",x"1e",
	x"10",x"0b",x"78",x"b1",x"20",x"d5",x"57",x"e1",x"c9",x"18",x"90",x"ed",x"73",x"3f",x"5c",x"fd",
	x"36",x"02",x"10",x"cd",x"af",x"0d",x"fd",x"cb",x"02",x"c6",x"fd",x"46",x"31",x"cd",x"44",x"0e",
	x"fd",x"cb",x"02",x"86",x"fd",x"cb",x"30",x"c6",x"2a",x"49",x"5c",x"ed",x"5b",x"6c",x"5c",x"a7",
	x"ed",x"52",x"19",x"38",x"22",x"d5",x"cd",x"6e",x"19",x"11",x"c0",x"02",x"eb",x"ed",x"52",x"e3",
	x"cd",x"6e",x"19",x"c1",x"c5",x"cd",x"b8",x"19",x"c1",x"09",x"38",x"0e",x"eb",x"56",x"23",x"5e",
	x"2b",x"ed",x"53",x"6c",x"5c",x"18",x"ed",x"22",x"6c",x"5c",x"2a",x"6c",x"5c",x"cd",x"6e",x"19",
	x"28",x"01",x"eb",x"cd",x"33",x"18",x"fd",x"cb",x"02",x"a6",x"c9",x"3e",x"03",x"18",x"02",x"3e",
	x"02",x"fd",x"36",x"02",x"00",x"cd",x"30",x"25",x"c4",x"01",x"16",x"df",x"cd",x"70",x"20",x"38",
	x"14",x"df",x"fe",x"3b",x"28",x"04",x"fe",x"2c",x"20",x"06",x"e7",x"cd",x"82",x"1c",x"18",x"08",
	x"cd",x"e6",x"1c",x"18",x"03",x"cd",x"de",x"1c",x"cd",x"ee",x"1b",x"cd",x"99",x"1e",x"78",x"e6",
	x"3f",x"67",x"69",x"22",x"49",x"5c",x"cd",x"6e",x"19",x"1e",x"01",x"cd",x"55",x"18",x"d7",x"fd",
	x"cb",x"02",x"66",x"28",x"f6",x"3a",x"6b",x"5c",x"fd",x"96",x"4f",x"20",x"ee",x"ab",x"c8",x"e5",
	x"d5",x"21",x"6c",x"5c",x"cd",x"0f",x"19",x"d1",x"e1",x"18",x"e0",x"ed",x"4b",x"49",x"5c",x"cd",
	x"80",x"19",x"16",x"3e",x"28",x"05",x"11",x"00",x"00",x"cb",x"13",x"fd",x"73",x"2d",x"7e",x"fe",
	x"40",x"c1",x"d0",x"c5",x"cd",x"28",x"1a",x"23",x"23",x"23",x"fd",x"cb",x"01",x"86",x"7a",x"a7",
	x"28",x"05",x"d7",x"fd",x"cb",x"01",x"c6",x"d5",x"eb",x"fd",x"cb",x"30",x"96",x"21",x"3b",x"5c",
	x"cb",x"96",x"fd",x"cb",x"37",x"6e",x"28",x"02",x"cb",x"d6",x"2a",x"5f",x"5c",x"a7",x"ed",x"52",
	x"20",x"05",x"3e",x"3f",x"cd",x"c1",x"18",x"cd",x"e1",x"18",x"eb",x"7e",x"cd",x"b6",x"18",x"23",
	x"fe",x"0d",x"28",x"06",x"eb",x"cd",x"37",x"19",x"18",x"e0",x"d1",x"c9",x"fe",x"0e",x"c0",x"23",
	x"23",x"23",x"23",x"23",x"23",x"7e",x"c9",x"d9",x"2a",x"8f",x"5c",x"e5",x"cb",x"bc",x"cb",x"fd",
	x"22",x"8f",x"5c",x"21",x"91",x"5c",x"56",x"d5",x"36",x"00",x"cd",x"f4",x"09",x"e1",x"fd",x"74",
	x"57",x"e1",x"22",x"8f",x"5c",x"d9",x"c9",x"2a",x"5b",x"5c",x"a7",x"ed",x"52",x"c0",x"3a",x"41",
	x"5c",x"cb",x"07",x"28",x"04",x"c6",x"43",x"18",x"16",x"21",x"3b",x"5c",x"cb",x"9e",x"3e",x"4b",
	x"cb",x"56",x"28",x"0b",x"cb",x"de",x"3c",x"fd",x"cb",x"30",x"5e",x"28",x"02",x"3e",x"43",x"d5",
	x"cd",x"c1",x"18",x"d1",x"c9",x"5e",x"23",x"56",x"e5",x"eb",x"23",x"cd",x"6e",x"19",x"cd",x"95",
	x"16",x"e1",x"fd",x"cb",x"37",x"6e",x"c0",x"72",x"2b",x"73",x"c9",x"7b",x"a7",x"f8",x"18",x"0d",
	x"af",x"09",x"3c",x"38",x"fc",x"ed",x"42",x"3d",x"28",x"f1",x"c3",x"ef",x"15",x"cd",x"1b",x"2d",
	x"30",x"30",x"fe",x"21",x"38",x"2c",x"fd",x"cb",x"01",x"96",x"fe",x"cb",x"28",x"24",x"fe",x"3a",
	x"20",x"0e",x"fd",x"cb",x"37",x"6e",x"20",x"16",x"fd",x"cb",x"30",x"56",x"28",x"14",x"18",x"0e",
	x"fe",x"22",x"20",x"0a",x"f5",x"3a",x"6a",x"5c",x"ee",x"04",x"32",x"6a",x"5c",x"f1",x"fd",x"cb",
	x"01",x"d6",x"d7",x"c9",x"e5",x"2a",x"53",x"5c",x"54",x"5d",x"c1",x"cd",x"80",x"19",x"d0",x"c5",
	x"cd",x"b8",x"19",x"eb",x"18",x"f4",x"7e",x"b8",x"c0",x"23",x"7e",x"2b",x"b9",x"c9",x"23",x"23",
	x"23",x"22",x"5d",x"5c",x"0e",x"00",x"15",x"c8",x"e7",x"bb",x"20",x"04",x"a7",x"c9",x"23",x"7e",
	x"cd",x"b6",x"18",x"22",x"5d",x"5c",x"fe",x"22",x"20",x"01",x"0d",x"fe",x"3a",x"28",x"04",x"fe",
	x"cb",x"20",x"04",x"cb",x"41",x"28",x"df",x"fe",x"0d",x"20",x"e3",x"15",x"37",x"c9",x"e5",x"7e",
	x"fe",x"40",x"38",x"17",x"cb",x"6f",x"28",x"14",x"87",x"fa",x"c7",x"19",x"3f",x"01",x"05",x"00",
	x"30",x"02",x"0e",x"12",x"17",x"23",x"7e",x"30",x"fb",x"18",x"06",x"23",x"23",x"4e",x"23",x"46",
	x"23",x"09",x"d1",x"a7",x"ed",x"52",x"44",x"4d",x"19",x"eb",x"c9",x"cd",x"dd",x"19",x"c5",x"78",
	x"2f",x"47",x"79",x"2f",x"4f",x"03",x"cd",x"64",x"16",x"eb",x"e1",x"19",x"d5",x"ed",x"b0",x"e1",
	x"c9",x"2a",x"59",x"5c",x"2b",x"22",x"5d",x"5c",x"e7",x"21",x"92",x"5c",x"22",x"65",x"5c",x"cd",
	x"3b",x"2d",x"cd",x"a2",x"2d",x"38",x"04",x"21",x"f0",x"d8",x"09",x"da",x"8a",x"1c",x"c3",x"c5",
	x"16",x"d5",x"e5",x"af",x"cb",x"78",x"20",x"20",x"60",x"69",x"1e",x"ff",x"18",x"08",x"d5",x"56",
	x"23",x"5e",x"e5",x"eb",x"1e",x"20",x"01",x"18",x"fc",x"cd",x"2a",x"19",x"01",x"9c",x"ff",x"cd",
	x"2a",x"19",x"0e",x"f6",x"cd",x"2a",x"19",x"7d",x"cd",x"ef",x"15",x"e1",x"d1",x"c9",x"b1",x"cb",
	x"bc",x"bf",x"c4",x"af",x"b4",x"93",x"91",x"92",x"95",x"98",x"98",x"98",x"98",x"98",x"98",x"98",
	x"7f",x"81",x"2e",x"6c",x"6e",x"70",x"48",x"94",x"56",x"3f",x"41",x"2b",x"17",x"1f",x"37",x"77",
	x"44",x"0f",x"59",x"2b",x"43",x"2d",x"51",x"3a",x"6d",x"42",x"0d",x"49",x"5c",x"44",x"15",x"5d",
	x"01",x"3d",x"02",x"06",x"00",x"67",x"1e",x"06",x"cb",x"05",x"f0",x"1c",x"06",x"00",x"ed",x"1e",
	x"00",x"ee",x"1c",x"00",x"23",x"1f",x"04",x"3d",x"06",x"cc",x"06",x"05",x"03",x"1d",x"04",x"00",
	x"ab",x"1d",x"05",x"cd",x"1f",x"05",x"89",x"20",x"05",x"02",x"2c",x"05",x"b2",x"1b",x"00",x"b7",
	x"11",x"03",x"a1",x"1e",x"05",x"f9",x"17",x"08",x"00",x"80",x"1e",x"03",x"4f",x"1e",x"00",x"5f",
	x"1e",x"03",x"ac",x"1e",x"00",x"6b",x"0d",x"09",x"00",x"dc",x"22",x"06",x"00",x"3a",x"1f",x"05",
	x"ed",x"1d",x"05",x"27",x"1e",x"03",x"42",x"1e",x"09",x"05",x"82",x"23",x"00",x"ac",x"0e",x"05",
	x"c9",x"1f",x"05",x"f5",x"17",x"0b",x"0b",x"0b",x"0b",x"08",x"00",x"f8",x"03",x"09",x"05",x"20",
	x"23",x"07",x"07",x"07",x"07",x"07",x"07",x"08",x"00",x"7a",x"1e",x"06",x"00",x"94",x"22",x"05",
	x"60",x"1f",x"06",x"2c",x"0a",x"00",x"36",x"17",x"06",x"00",x"e5",x"16",x"0a",x"00",x"93",x"17",
	x"0a",x"2c",x"0a",x"00",x"93",x"17",x"0a",x"00",x"93",x"17",x"00",x"93",x"17",x"fd",x"cb",x"01",
	x"be",x"cd",x"fb",x"19",x"af",x"32",x"47",x"5c",x"3d",x"32",x"3a",x"5c",x"18",x"01",x"e7",x"cd",
	x"bf",x"16",x"fd",x"34",x"0d",x"fa",x"8a",x"1c",x"df",x"06",x"00",x"fe",x"0d",x"28",x"7a",x"fe",
	x"3a",x"28",x"eb",x"21",x"76",x"1b",x"e5",x"4f",x"e7",x"79",x"d6",x"ce",x"da",x"8a",x"1c",x"4f",
	x"21",x"48",x"1a",x"09",x"4e",x"09",x"18",x"03",x"2a",x"74",x"5c",x"7e",x"23",x"22",x"74",x"5c",
	x"01",x"52",x"1b",x"c5",x"4f",x"fe",x"20",x"30",x"0c",x"21",x"01",x"1c",x"06",x"00",x"09",x"4e",
	x"09",x"e5",x"df",x"05",x"c9",x"df",x"b9",x"c2",x"8a",x"1c",x"e7",x"c9",x"cd",x"54",x"1f",x"38",
	x"02",x"cf",x"14",x"fd",x"cb",x"0a",x"7e",x"20",x"71",x"2a",x"42",x"5c",x"cb",x"7c",x"28",x"14",
	x"21",x"fe",x"ff",x"22",x"45",x"5c",x"2a",x"61",x"5c",x"2b",x"ed",x"5b",x"59",x"5c",x"1b",x"3a",
	x"44",x"5c",x"18",x"33",x"cd",x"6e",x"19",x"3a",x"44",x"5c",x"28",x"19",x"a7",x"20",x"43",x"47",
	x"7e",x"e6",x"c0",x"78",x"28",x"0f",x"cf",x"ff",x"c1",x"cd",x"30",x"25",x"c8",x"2a",x"55",x"5c",
	x"3e",x"c0",x"a6",x"c0",x"af",x"fe",x"01",x"ce",x"00",x"56",x"23",x"5e",x"ed",x"53",x"45",x"5c",
	x"23",x"5e",x"23",x"56",x"eb",x"19",x"23",x"22",x"55",x"5c",x"eb",x"22",x"5d",x"5c",x"57",x"1e",
	x"00",x"fd",x"36",x"0a",x"ff",x"15",x"fd",x"72",x"0d",x"ca",x"28",x"1b",x"14",x"cd",x"8b",x"19",
	x"28",x"08",x"cf",x"16",x"cd",x"30",x"25",x"c0",x"c1",x"c1",x"df",x"fe",x"0d",x"28",x"ba",x"fe",
	x"3a",x"ca",x"28",x"1b",x"c3",x"8a",x"1c",x"0f",x"1d",x"4b",x"09",x"67",x"0b",x"7b",x"8e",x"71",
	x"b4",x"81",x"cf",x"cd",x"de",x"1c",x"bf",x"c1",x"cc",x"ee",x"1b",x"eb",x"2a",x"74",x"5c",x"4e",
	x"23",x"46",x"eb",x"c5",x"c9",x"cd",x"b2",x"28",x"fd",x"36",x"37",x"00",x"30",x"08",x"fd",x"cb",
	x"37",x"ce",x"20",x"18",x"cf",x"01",x"cc",x"96",x"29",x"fd",x"cb",x"01",x"76",x"20",x"0d",x"af",
	x"cd",x"30",x"25",x"c4",x"f1",x"2b",x"21",x"71",x"5c",x"b6",x"77",x"eb",x"ed",x"43",x"72",x"5c",
	x"22",x"4d",x"5c",x"c9",x"c1",x"cd",x"56",x"1c",x"cd",x"ee",x"1b",x"c9",x"3a",x"3b",x"5c",x"f5",
	x"cd",x"fb",x"24",x"f1",x"fd",x"56",x"01",x"aa",x"e6",x"40",x"20",x"24",x"cb",x"7a",x"c2",x"ff",
	x"2a",x"c9",x"cd",x"b2",x"28",x"f5",x"79",x"f6",x"9f",x"3c",x"20",x"14",x"f1",x"18",x"a9",x"e7",
	x"cd",x"82",x"1c",x"fe",x"2c",x"20",x"09",x"e7",x"cd",x"fb",x"24",x"fd",x"cb",x"01",x"76",x"c0",
	x"cf",x"0b",x"cd",x"fb",x"24",x"fd",x"cb",x"01",x"76",x"c8",x"18",x"f4",x"fd",x"cb",x"01",x"7e",
	x"fd",x"cb",x"02",x"86",x"c4",x"4d",x"0d",x"f1",x"3a",x"74",x"5c",x"d6",x"13",x"cd",x"fc",x"21",
	x"cd",x"ee",x"1b",x"2a",x"8f",x"5c",x"22",x"8d",x"5c",x"21",x"91",x"5c",x"7e",x"07",x"ae",x"e6",
	x"aa",x"ae",x"77",x"c9",x"cd",x"30",x"25",x"28",x"13",x"fd",x"cb",x"02",x"86",x"cd",x"4d",x"0d",
	x"21",x"90",x"5c",x"7e",x"f6",x"f8",x"77",x"fd",x"cb",x"57",x"b6",x"df",x"cd",x"e2",x"21",x"18",
	x"9f",x"c3",x"05",x"06",x"fe",x"0d",x"28",x"04",x"fe",x"3a",x"20",x"9c",x"cd",x"30",x"25",x"c8",
	x"ef",x"a0",x"38",x"c9",x"cf",x"08",x"c1",x"cd",x"30",x"25",x"28",x"0a",x"ef",x"02",x"38",x"eb",
	x"cd",x"e9",x"34",x"da",x"b3",x"1b",x"c3",x"29",x"1b",x"fe",x"cd",x"20",x"09",x"e7",x"cd",x"82",
	x"1c",x"cd",x"ee",x"1b",x"18",x"06",x"cd",x"ee",x"1b",x"ef",x"a1",x"38",x"ef",x"c0",x"02",x"01",
	x"e0",x"01",x"38",x"cd",x"ff",x"2a",x"22",x"68",x"5c",x"2b",x"7e",x"cb",x"fe",x"01",x"06",x"00",
	x"09",x"07",x"38",x"06",x"0e",x"0d",x"cd",x"55",x"16",x"23",x"e5",x"ef",x"02",x"02",x"38",x"e1",
	x"eb",x"0e",x"0a",x"ed",x"b0",x"2a",x"45",x"5c",x"eb",x"73",x"23",x"72",x"fd",x"56",x"0d",x"14",
	x"23",x"72",x"cd",x"da",x"1d",x"d0",x"fd",x"46",x"38",x"2a",x"45",x"5c",x"22",x"42",x"5c",x"3a",
	x"47",x"5c",x"ed",x"44",x"57",x"2a",x"5d",x"5c",x"1e",x"f3",x"c5",x"ed",x"4b",x"55",x"5c",x"cd",
	x"86",x"1d",x"ed",x"43",x"55",x"5c",x"c1",x"38",x"11",x"e7",x"f6",x"20",x"b8",x"28",x"03",x"e7",
	x"18",x"e8",x"e7",x"3e",x"01",x"92",x"32",x"44",x"5c",x"c9",x"cf",x"11",x"7e",x"fe",x"3a",x"28",
	x"18",x"23",x"7e",x"e6",x"c0",x"37",x"c0",x"46",x"23",x"4e",x"ed",x"43",x"42",x"5c",x"23",x"4e",
	x"23",x"46",x"e5",x"09",x"44",x"4d",x"e1",x"16",x"00",x"c5",x"cd",x"8b",x"19",x"c1",x"d0",x"18",
	x"e0",x"fd",x"cb",x"37",x"4e",x"c2",x"2e",x"1c",x"2a",x"4d",x"5c",x"cb",x"7e",x"28",x"1f",x"23",
	x"22",x"68",x"5c",x"ef",x"e0",x"e2",x"0f",x"c0",x"02",x"38",x"cd",x"da",x"1d",x"d8",x"2a",x"68",
	x"5c",x"11",x"0f",x"00",x"19",x"5e",x"23",x"56",x"23",x"66",x"eb",x"c3",x"73",x"1e",x"cf",x"00",
	x"ef",x"e1",x"e0",x"e2",x"36",x"00",x"02",x"01",x"03",x"37",x"00",x"04",x"38",x"a7",x"c9",x"38",
	x"37",x"c9",x"e7",x"cd",x"1f",x"1c",x"cd",x"30",x"25",x"28",x"29",x"df",x"22",x"5f",x"5c",x"2a",
	x"57",x"5c",x"7e",x"fe",x"2c",x"28",x"09",x"1e",x"e4",x"cd",x"86",x"1d",x"30",x"02",x"cf",x"0d",
	x"cd",x"77",x"00",x"cd",x"56",x"1c",x"df",x"22",x"57",x"5c",x"2a",x"5f",x"5c",x"fd",x"36",x"26",
	x"00",x"cd",x"78",x"00",x"df",x"fe",x"2c",x"28",x"c9",x"cd",x"ee",x"1b",x"c9",x"cd",x"30",x"25",
	x"20",x"0b",x"cd",x"fb",x"24",x"fe",x"2c",x"c4",x"ee",x"1b",x"e7",x"18",x"f5",x"3e",x"e4",x"47",
	x"ed",x"b9",x"11",x"00",x"02",x"c3",x"8b",x"19",x"cd",x"99",x"1e",x"60",x"69",x"cd",x"6e",x"19",
	x"2b",x"22",x"57",x"5c",x"c9",x"cd",x"99",x"1e",x"78",x"b1",x"20",x"04",x"ed",x"4b",x"78",x"5c",
	x"ed",x"43",x"76",x"5c",x"c9",x"2a",x"6e",x"5c",x"fd",x"56",x"36",x"18",x"0c",x"cd",x"99",x"1e",
	x"60",x"69",x"16",x"00",x"7c",x"fe",x"f0",x"30",x"2c",x"22",x"42",x"5c",x"fd",x"72",x"0a",x"c9",
	x"cd",x"85",x"1e",x"ed",x"79",x"c9",x"cd",x"85",x"1e",x"02",x"c9",x"cd",x"d5",x"2d",x"38",x"15",
	x"28",x"02",x"ed",x"44",x"f5",x"cd",x"99",x"1e",x"f1",x"c9",x"cd",x"d5",x"2d",x"18",x"03",x"cd",
	x"a2",x"2d",x"38",x"01",x"c8",x"cf",x"0a",x"cd",x"67",x"1e",x"01",x"00",x"00",x"cd",x"45",x"1e",
	x"18",x"03",x"cd",x"99",x"1e",x"78",x"b1",x"20",x"04",x"ed",x"4b",x"b2",x"5c",x"c5",x"ed",x"5b",
	x"4b",x"5c",x"2a",x"59",x"5c",x"2b",x"cd",x"e5",x"19",x"cd",x"6b",x"0d",x"2a",x"65",x"5c",x"11",
	x"32",x"00",x"19",x"d1",x"ed",x"52",x"30",x"08",x"2a",x"b4",x"5c",x"a7",x"ed",x"52",x"30",x"02",
	x"cf",x"15",x"eb",x"22",x"b2",x"5c",x"d1",x"c1",x"36",x"3e",x"2b",x"f9",x"c5",x"ed",x"73",x"3d",
	x"5c",x"eb",x"e9",x"d1",x"fd",x"66",x"0d",x"24",x"e3",x"33",x"ed",x"4b",x"45",x"5c",x"c5",x"e5",
	x"ed",x"73",x"3d",x"5c",x"d5",x"cd",x"67",x"1e",x"01",x"14",x"00",x"2a",x"65",x"5c",x"09",x"38",
	x"0a",x"eb",x"21",x"50",x"00",x"19",x"38",x"03",x"ed",x"72",x"d8",x"2e",x"03",x"c3",x"55",x"00",
	x"01",x"00",x"00",x"cd",x"05",x"1f",x"44",x"4d",x"c9",x"c1",x"e1",x"d1",x"7a",x"fe",x"3e",x"28",
	x"0b",x"3b",x"e3",x"eb",x"ed",x"73",x"3d",x"5c",x"c5",x"c3",x"73",x"1e",x"d5",x"e5",x"cf",x"06",
	x"cd",x"99",x"1e",x"76",x"0b",x"78",x"b1",x"28",x"0c",x"78",x"a1",x"3c",x"20",x"01",x"03",x"fd",
	x"cb",x"01",x"6e",x"28",x"ee",x"fd",x"cb",x"01",x"ae",x"c9",x"3e",x"7f",x"db",x"fe",x"1f",x"d8",
	x"3e",x"fe",x"db",x"fe",x"1f",x"c9",x"cd",x"30",x"25",x"28",x"05",x"3e",x"ce",x"c3",x"39",x"1e",
	x"fd",x"cb",x"01",x"f6",x"cd",x"8d",x"2c",x"30",x"16",x"e7",x"fe",x"24",x"20",x"05",x"fd",x"cb",
	x"01",x"b6",x"e7",x"fe",x"28",x"20",x"3c",x"e7",x"fe",x"29",x"28",x"20",x"cd",x"8d",x"2c",x"d2",
	x"8a",x"1c",x"eb",x"e7",x"fe",x"24",x"20",x"02",x"eb",x"e7",x"eb",x"01",x"06",x"00",x"cd",x"55",
	x"16",x"23",x"23",x"36",x"0e",x"fe",x"2c",x"20",x"03",x"e7",x"18",x"e0",x"fe",x"29",x"20",x"13",
	x"e7",x"fe",x"3d",x"20",x"0e",x"e7",x"3a",x"3b",x"5c",x"f5",x"cd",x"fb",x"24",x"f1",x"fd",x"ae",
	x"01",x"e6",x"40",x"c2",x"8a",x"1c",x"cd",x"ee",x"1b",x"cd",x"30",x"25",x"e1",x"c8",x"e9",x"3e",
	x"03",x"18",x"02",x"3e",x"02",x"cd",x"30",x"25",x"c4",x"01",x"16",x"cd",x"4d",x"0d",x"cd",x"df",
	x"1f",x"cd",x"ee",x"1b",x"c9",x"df",x"cd",x"45",x"20",x"28",x"0d",x"cd",x"4e",x"20",x"28",x"fb",
	x"cd",x"fc",x"1f",x"cd",x"4e",x"20",x"28",x"f3",x"fe",x"29",x"c8",x"cd",x"c3",x"1f",x"3e",x"0d",
	x"d7",x"c9",x"df",x"fe",x"ac",x"20",x"0d",x"cd",x"79",x"1c",x"cd",x"c3",x"1f",x"cd",x"07",x"23",
	x"3e",x"16",x"18",x"10",x"fe",x"ad",x"20",x"12",x"e7",x"cd",x"82",x"1c",x"cd",x"c3",x"1f",x"cd",
	x"99",x"1e",x"3e",x"17",x"d7",x"79",x"d7",x"78",x"d7",x"c9",x"cd",x"f2",x"21",x"d0",x"cd",x"70",
	x"20",x"d0",x"cd",x"fb",x"24",x"cd",x"c3",x"1f",x"fd",x"cb",x"01",x"76",x"cc",x"f1",x"2b",x"c2",
	x"e3",x"2d",x"78",x"b1",x"0b",x"c8",x"1a",x"13",x"d7",x"18",x"f7",x"fe",x"29",x"c8",x"fe",x"0d",
	x"c8",x"fe",x"3a",x"c9",x"df",x"fe",x"3b",x"28",x"14",x"fe",x"2c",x"20",x"0a",x"cd",x"30",x"25",
	x"28",x"0b",x"3e",x"06",x"d7",x"18",x"06",x"fe",x"27",x"c0",x"cd",x"f5",x"1f",x"e7",x"cd",x"45",
	x"20",x"20",x"01",x"c1",x"bf",x"c9",x"fe",x"23",x"37",x"c0",x"e7",x"cd",x"82",x"1c",x"a7",x"cd",
	x"c3",x"1f",x"cd",x"94",x"1e",x"fe",x"10",x"d2",x"0e",x"16",x"cd",x"01",x"16",x"a7",x"c9",x"cd",
	x"30",x"25",x"28",x"08",x"3e",x"01",x"cd",x"01",x"16",x"cd",x"6e",x"0d",x"fd",x"36",x"02",x"01",
	x"cd",x"c1",x"20",x"cd",x"ee",x"1b",x"ed",x"4b",x"88",x"5c",x"3a",x"6b",x"5c",x"b8",x"38",x"03",
	x"0e",x"21",x"47",x"ed",x"43",x"88",x"5c",x"3e",x"19",x"90",x"32",x"8c",x"5c",x"fd",x"cb",x"02",
	x"86",x"cd",x"d9",x"0d",x"c3",x"6e",x"0d",x"cd",x"4e",x"20",x"28",x"fb",x"fe",x"28",x"20",x"0e",
	x"e7",x"cd",x"df",x"1f",x"df",x"fe",x"29",x"c2",x"8a",x"1c",x"e7",x"c3",x"b2",x"21",x"fe",x"ca",
	x"20",x"11",x"e7",x"cd",x"1f",x"1c",x"fd",x"cb",x"37",x"fe",x"fd",x"cb",x"01",x"76",x"c2",x"8a",
	x"1c",x"18",x"0d",x"cd",x"8d",x"2c",x"d2",x"af",x"21",x"cd",x"1f",x"1c",x"fd",x"cb",x"37",x"be",
	x"cd",x"30",x"25",x"ca",x"b2",x"21",x"cd",x"bf",x"16",x"21",x"71",x"5c",x"cb",x"b6",x"cb",x"ee",
	x"01",x"01",x"00",x"cb",x"7e",x"20",x"0b",x"3a",x"3b",x"5c",x"e6",x"40",x"20",x"02",x"0e",x"03",
	x"b6",x"77",x"f7",x"36",x"0d",x"79",x"0f",x"0f",x"30",x"05",x"3e",x"22",x"12",x"2b",x"77",x"22",
	x"5b",x"5c",x"fd",x"cb",x"37",x"7e",x"20",x"2c",x"2a",x"5d",x"5c",x"e5",x"2a",x"3d",x"5c",x"e5",
	x"21",x"3a",x"21",x"e5",x"fd",x"cb",x"30",x"66",x"28",x"04",x"ed",x"73",x"3d",x"5c",x"2a",x"61",
	x"5c",x"cd",x"a7",x"11",x"fd",x"36",x"00",x"ff",x"cd",x"2c",x"0f",x"fd",x"cb",x"01",x"be",x"cd",
	x"b9",x"21",x"18",x"03",x"cd",x"2c",x"0f",x"fd",x"36",x"22",x"00",x"cd",x"d6",x"21",x"20",x"0a",
	x"cd",x"1d",x"11",x"ed",x"4b",x"82",x"5c",x"cd",x"d9",x"0d",x"21",x"71",x"5c",x"cb",x"ae",x"cb",
	x"7e",x"cb",x"be",x"20",x"1c",x"e1",x"e1",x"22",x"3d",x"5c",x"e1",x"22",x"5f",x"5c",x"fd",x"cb",
	x"01",x"fe",x"cd",x"b9",x"21",x"2a",x"5f",x"5c",x"fd",x"36",x"26",x"00",x"22",x"5d",x"5c",x"18",
	x"17",x"2a",x"63",x"5c",x"ed",x"5b",x"61",x"5c",x"37",x"ed",x"52",x"44",x"4d",x"cd",x"b2",x"2a",
	x"cd",x"ff",x"2a",x"18",x"03",x"cd",x"fc",x"1f",x"cd",x"4e",x"20",x"ca",x"c1",x"20",x"c9",x"2a",
	x"61",x"5c",x"22",x"5d",x"5c",x"df",x"fe",x"e2",x"28",x"0c",x"3a",x"71",x"5c",x"cd",x"59",x"1c",
	x"df",x"fe",x"0d",x"c8",x"cf",x"0b",x"cd",x"30",x"25",x"c8",x"cf",x"10",x"2a",x"51",x"5c",x"23",
	x"23",x"23",x"23",x"7e",x"fe",x"4b",x"c9",x"e7",x"cd",x"f2",x"21",x"d8",x"df",x"fe",x"2c",x"28",
	x"f6",x"fe",x"3b",x"28",x"f2",x"c3",x"8a",x"1c",x"fe",x"d9",x"d8",x"fe",x"df",x"3f",x"d8",x"f5",
	x"e7",x"f1",x"d6",x"c9",x"f5",x"cd",x"82",x"1c",x"f1",x"a7",x"cd",x"c3",x"1f",x"f5",x"cd",x"94",
	x"1e",x"57",x"f1",x"d7",x"7a",x"d7",x"c9",x"d6",x"11",x"ce",x"00",x"28",x"1d",x"d6",x"02",x"ce",
	x"00",x"28",x"56",x"fe",x"01",x"7a",x"06",x"01",x"20",x"04",x"07",x"07",x"06",x"04",x"4f",x"7a",
	x"fe",x"02",x"30",x"16",x"79",x"21",x"91",x"5c",x"18",x"38",x"7a",x"06",x"07",x"38",x"05",x"07",
	x"07",x"07",x"06",x"38",x"4f",x"7a",x"fe",x"0a",x"38",x"02",x"cf",x"13",x"21",x"8f",x"5c",x"fe",
	x"08",x"38",x"0b",x"7e",x"28",x"07",x"b0",x"2f",x"e6",x"24",x"28",x"01",x"78",x"4f",x"79",x"cd",
	x"6c",x"22",x"3e",x"07",x"ba",x"9f",x"cd",x"6c",x"22",x"07",x"07",x"e6",x"50",x"47",x"3e",x"08",
	x"ba",x"9f",x"ae",x"a0",x"ae",x"77",x"23",x"78",x"c9",x"9f",x"7a",x"0f",x"06",x"80",x"20",x"03",
	x"0f",x"06",x"40",x"4f",x"7a",x"fe",x"08",x"28",x"04",x"fe",x"02",x"30",x"bd",x"79",x"21",x"8f",
	x"5c",x"cd",x"6c",x"22",x"79",x"0f",x"0f",x"0f",x"18",x"d8",x"cd",x"94",x"1e",x"fe",x"08",x"30",
	x"a9",x"d3",x"fe",x"07",x"07",x"07",x"cb",x"6f",x"20",x"02",x"ee",x"07",x"32",x"48",x"5c",x"c9",
	x"3e",x"af",x"90",x"da",x"f9",x"24",x"47",x"a7",x"1f",x"37",x"1f",x"a7",x"1f",x"a8",x"e6",x"f8",
	x"a8",x"67",x"79",x"07",x"07",x"07",x"a8",x"e6",x"c7",x"a8",x"07",x"07",x"6f",x"79",x"e6",x"07",
	x"c9",x"cd",x"07",x"23",x"cd",x"aa",x"22",x"47",x"04",x"7e",x"07",x"10",x"fd",x"e6",x"01",x"c3",
	x"28",x"2d",x"cd",x"07",x"23",x"cd",x"e5",x"22",x"c3",x"4d",x"0d",x"ed",x"43",x"7d",x"5c",x"cd",
	x"aa",x"22",x"47",x"04",x"3e",x"fe",x"0f",x"10",x"fd",x"47",x"7e",x"fd",x"4e",x"57",x"cb",x"41",
	x"20",x"01",x"a0",x"cb",x"51",x"20",x"02",x"a8",x"2f",x"77",x"c3",x"db",x"0b",x"cd",x"14",x"23",
	x"47",x"c5",x"cd",x"14",x"23",x"59",x"c1",x"51",x"4f",x"c9",x"cd",x"d5",x"2d",x"da",x"f9",x"24",
	x"0e",x"01",x"c8",x"0e",x"ff",x"c9",x"df",x"fe",x"2c",x"c2",x"8a",x"1c",x"e7",x"cd",x"82",x"1c",
	x"cd",x"ee",x"1b",x"ef",x"2a",x"3d",x"38",x"7e",x"fe",x"81",x"30",x"05",x"ef",x"02",x"38",x"18",
	x"a1",x"ef",x"a3",x"38",x"36",x"83",x"ef",x"c5",x"02",x"38",x"cd",x"7d",x"24",x"c5",x"ef",x"31",
	x"e1",x"04",x"38",x"7e",x"fe",x"80",x"30",x"08",x"ef",x"02",x"02",x"38",x"c1",x"c3",x"dc",x"22",
	x"ef",x"c2",x"01",x"c0",x"02",x"03",x"01",x"e0",x"0f",x"c0",x"01",x"31",x"e0",x"01",x"31",x"e0",
	x"a0",x"c1",x"02",x"38",x"fd",x"34",x"62",x"cd",x"94",x"1e",x"6f",x"e5",x"cd",x"94",x"1e",x"e1",
	x"67",x"22",x"7d",x"5c",x"c1",x"c3",x"20",x"24",x"df",x"fe",x"2c",x"28",x"06",x"cd",x"ee",x"1b",
	x"c3",x"77",x"24",x"e7",x"cd",x"82",x"1c",x"cd",x"ee",x"1b",x"ef",x"c5",x"a2",x"04",x"1f",x"31",
	x"30",x"30",x"00",x"06",x"02",x"38",x"c3",x"77",x"24",x"c0",x"02",x"c1",x"02",x"31",x"2a",x"e1",
	x"01",x"e1",x"2a",x"0f",x"e0",x"05",x"2a",x"e0",x"01",x"3d",x"38",x"7e",x"fe",x"81",x"30",x"07",
	x"ef",x"02",x"02",x"38",x"c3",x"77",x"24",x"cd",x"7d",x"24",x"c5",x"ef",x"02",x"e1",x"01",x"05",
	x"c1",x"02",x"01",x"31",x"e1",x"04",x"c2",x"02",x"01",x"31",x"e1",x"04",x"e2",x"e5",x"e0",x"03",
	x"a2",x"04",x"31",x"1f",x"c5",x"02",x"20",x"c0",x"02",x"c2",x"02",x"c1",x"e5",x"04",x"e0",x"e2",
	x"04",x"0f",x"e1",x"01",x"c1",x"02",x"e0",x"04",x"e2",x"e5",x"04",x"03",x"c2",x"2a",x"e1",x"2a",
	x"0f",x"02",x"38",x"1a",x"fe",x"81",x"c1",x"da",x"77",x"24",x"c5",x"ef",x"01",x"38",x"3a",x"7d",
	x"5c",x"cd",x"28",x"2d",x"ef",x"c0",x"0f",x"01",x"38",x"3a",x"7e",x"5c",x"cd",x"28",x"2d",x"ef",
	x"c5",x"0f",x"e0",x"e5",x"38",x"c1",x"05",x"28",x"3c",x"18",x"14",x"ef",x"e1",x"31",x"e3",x"04",
	x"e2",x"e4",x"04",x"03",x"c1",x"02",x"e4",x"04",x"e2",x"e3",x"04",x"0f",x"c2",x"02",x"38",x"c5",
	x"ef",x"c0",x"02",x"e1",x"0f",x"31",x"38",x"3a",x"7d",x"5c",x"cd",x"28",x"2d",x"ef",x"03",x"e0",
	x"e2",x"0f",x"c0",x"01",x"e0",x"38",x"3a",x"7e",x"5c",x"cd",x"28",x"2d",x"ef",x"03",x"38",x"cd",
	x"b7",x"24",x"c1",x"10",x"c6",x"ef",x"02",x"02",x"01",x"38",x"3a",x"7d",x"5c",x"cd",x"28",x"2d",
	x"ef",x"03",x"01",x"38",x"3a",x"7e",x"5c",x"cd",x"28",x"2d",x"ef",x"03",x"38",x"cd",x"b7",x"24",
	x"c3",x"4d",x"0d",x"ef",x"31",x"28",x"34",x"32",x"00",x"01",x"05",x"e5",x"01",x"05",x"2a",x"38",
	x"cd",x"d5",x"2d",x"38",x"06",x"e6",x"fc",x"c6",x"04",x"30",x"02",x"3e",x"fc",x"f5",x"cd",x"28",
	x"2d",x"ef",x"e5",x"01",x"05",x"31",x"1f",x"c4",x"02",x"31",x"a2",x"04",x"1f",x"c1",x"01",x"c0",
	x"02",x"31",x"04",x"31",x"0f",x"a1",x"03",x"1b",x"c3",x"02",x"38",x"c1",x"c9",x"cd",x"07",x"23",
	x"79",x"b8",x"30",x"06",x"69",x"d5",x"af",x"5f",x"18",x"07",x"b1",x"c8",x"68",x"41",x"d5",x"16",
	x"00",x"60",x"78",x"1f",x"85",x"38",x"03",x"bc",x"38",x"07",x"94",x"4f",x"d9",x"c1",x"c5",x"18",
	x"04",x"4f",x"d5",x"d9",x"c1",x"2a",x"7d",x"5c",x"78",x"84",x"47",x"79",x"3c",x"85",x"38",x"0d",
	x"28",x"0d",x"3d",x"4f",x"cd",x"e5",x"22",x"d9",x"79",x"10",x"d9",x"d1",x"c9",x"28",x"f3",x"cf",
	x"0a",x"df",x"06",x"00",x"c5",x"4f",x"21",x"96",x"25",x"cd",x"dc",x"16",x"79",x"d2",x"84",x"26",
	x"06",x"00",x"4e",x"09",x"e9",x"cd",x"74",x"00",x"03",x"fe",x"0d",x"ca",x"8a",x"1c",x"fe",x"22",
	x"20",x"f3",x"cd",x"74",x"00",x"fe",x"22",x"c9",x"e7",x"fe",x"28",x"20",x"06",x"cd",x"79",x"1c",
	x"df",x"fe",x"29",x"c2",x"8a",x"1c",x"fd",x"cb",x"01",x"7e",x"c9",x"cd",x"07",x"23",x"2a",x"36",
	x"5c",x"11",x"00",x"01",x"19",x"79",x"0f",x"0f",x"0f",x"e6",x"e0",x"a8",x"5f",x"79",x"e6",x"18",
	x"ee",x"40",x"57",x"06",x"60",x"c5",x"d5",x"e5",x"1a",x"ae",x"28",x"04",x"3c",x"20",x"1a",x"3d",
	x"4f",x"06",x"07",x"14",x"23",x"1a",x"ae",x"a9",x"20",x"0f",x"10",x"f7",x"c1",x"c1",x"c1",x"3e",
	x"80",x"90",x"01",x"01",x"00",x"f7",x"12",x"18",x"0a",x"e1",x"11",x"08",x"00",x"19",x"d1",x"c1",
	x"10",x"d3",x"48",x"c3",x"b2",x"2a",x"cd",x"07",x"23",x"79",x"0f",x"0f",x"0f",x"4f",x"e6",x"e0",
	x"a8",x"6f",x"79",x"e6",x"03",x"ee",x"58",x"67",x"7e",x"c3",x"28",x"2d",x"22",x"1c",x"28",x"4f",
	x"2e",x"f2",x"2b",x"12",x"a8",x"56",x"a5",x"57",x"a7",x"84",x"a6",x"8f",x"c4",x"e6",x"aa",x"bf",
	x"ab",x"c7",x"a9",x"ce",x"00",x"e7",x"c3",x"ff",x"24",x"df",x"23",x"e5",x"01",x"00",x"00",x"cd",
	x"0f",x"25",x"20",x"1b",x"cd",x"0f",x"25",x"28",x"fb",x"cd",x"30",x"25",x"28",x"11",x"f7",x"e1",
	x"d5",x"7e",x"23",x"12",x"13",x"fe",x"22",x"20",x"f8",x"7e",x"23",x"fe",x"22",x"28",x"f2",x"0b",
	x"d1",x"21",x"3b",x"5c",x"cb",x"b6",x"cb",x"7e",x"c4",x"b2",x"2a",x"c3",x"12",x"27",x"e7",x"cd",
	x"fb",x"24",x"fe",x"29",x"c2",x"8a",x"1c",x"e7",x"c3",x"12",x"27",x"c3",x"bd",x"27",x"cd",x"30",
	x"25",x"28",x"28",x"ed",x"4b",x"76",x"5c",x"cd",x"2b",x"2d",x"ef",x"a1",x"0f",x"34",x"37",x"16",
	x"04",x"34",x"80",x"41",x"00",x"00",x"80",x"32",x"02",x"a1",x"03",x"31",x"38",x"cd",x"a2",x"2d",
	x"ed",x"43",x"76",x"5c",x"7e",x"a7",x"28",x"03",x"d6",x"10",x"77",x"18",x"09",x"cd",x"30",x"25",
	x"28",x"04",x"ef",x"a3",x"38",x"34",x"e7",x"c3",x"c3",x"26",x"01",x"5a",x"10",x"e7",x"fe",x"23",
	x"ca",x"0d",x"27",x"21",x"3b",x"5c",x"cb",x"b6",x"cb",x"7e",x"28",x"1f",x"cd",x"8e",x"02",x"0e",
	x"00",x"20",x"13",x"cd",x"1e",x"03",x"30",x"0e",x"15",x"5f",x"cd",x"33",x"03",x"f5",x"01",x"01",
	x"00",x"f7",x"f1",x"12",x"0e",x"01",x"06",x"00",x"cd",x"b2",x"2a",x"c3",x"12",x"27",x"cd",x"22",
	x"25",x"c4",x"35",x"25",x"e7",x"c3",x"db",x"25",x"cd",x"22",x"25",x"c4",x"80",x"25",x"e7",x"18",
	x"48",x"cd",x"22",x"25",x"c4",x"cb",x"22",x"e7",x"18",x"3f",x"cd",x"88",x"2c",x"30",x"56",x"fe",
	x"41",x"30",x"3c",x"cd",x"30",x"25",x"20",x"23",x"cd",x"9b",x"2c",x"df",x"01",x"06",x"00",x"cd",
	x"55",x"16",x"23",x"36",x"0e",x"23",x"eb",x"2a",x"65",x"5c",x"0e",x"05",x"a7",x"ed",x"42",x"22",
	x"65",x"5c",x"ed",x"b0",x"eb",x"2b",x"cd",x"77",x"00",x"18",x"0e",x"df",x"23",x"7e",x"fe",x"0e",
	x"20",x"fa",x"23",x"cd",x"b4",x"33",x"22",x"5d",x"5c",x"fd",x"cb",x"01",x"f6",x"18",x"14",x"cd",
	x"b2",x"28",x"da",x"2e",x"1c",x"cc",x"96",x"29",x"3a",x"3b",x"5c",x"fe",x"c0",x"38",x"04",x"23",
	x"cd",x"b4",x"33",x"18",x"33",x"01",x"db",x"09",x"fe",x"2d",x"28",x"27",x"01",x"18",x"10",x"fe",
	x"ae",x"28",x"20",x"d6",x"af",x"da",x"8a",x"1c",x"01",x"f0",x"04",x"fe",x"14",x"28",x"14",x"d2",
	x"8a",x"1c",x"06",x"10",x"c6",x"dc",x"4f",x"fe",x"df",x"30",x"02",x"cb",x"b1",x"fe",x"ee",x"38",
	x"02",x"cb",x"b9",x"c5",x"e7",x"c3",x"ff",x"24",x"df",x"fe",x"28",x"20",x"0c",x"fd",x"cb",x"01",
	x"76",x"20",x"17",x"cd",x"52",x"2a",x"e7",x"18",x"f0",x"06",x"00",x"4f",x"21",x"95",x"27",x"cd",
	x"dc",x"16",x"30",x"06",x"4e",x"21",x"ed",x"26",x"09",x"46",x"d1",x"7a",x"b8",x"38",x"3a",x"a7",
	x"ca",x"18",x"00",x"c5",x"21",x"3b",x"5c",x"7b",x"fe",x"ed",x"20",x"06",x"cb",x"76",x"20",x"02",
	x"1e",x"99",x"d5",x"cd",x"30",x"25",x"28",x"09",x"7b",x"e6",x"3f",x"47",x"ef",x"3b",x"38",x"18",
	x"09",x"7b",x"fd",x"ae",x"01",x"e6",x"40",x"c2",x"8a",x"1c",x"d1",x"21",x"3b",x"5c",x"cb",x"f6",
	x"cb",x"7b",x"20",x"02",x"cb",x"b6",x"c1",x"18",x"c1",x"d5",x"79",x"fd",x"cb",x"01",x"76",x"20",
	x"15",x"e6",x"3f",x"c6",x"08",x"4f",x"fe",x"10",x"20",x"04",x"cb",x"f1",x"18",x"08",x"38",x"d7",
	x"fe",x"17",x"28",x"02",x"cb",x"f9",x"c5",x"e7",x"c3",x"ff",x"24",x"2b",x"cf",x"2d",x"c3",x"2a",
	x"c4",x"2f",x"c5",x"5e",x"c6",x"3d",x"ce",x"3e",x"cc",x"3c",x"cd",x"c7",x"c9",x"c8",x"ca",x"c9",
	x"cb",x"c5",x"c7",x"c6",x"c8",x"00",x"06",x"08",x"08",x"0a",x"02",x"03",x"05",x"05",x"05",x"05",
	x"05",x"05",x"06",x"cd",x"30",x"25",x"20",x"35",x"e7",x"cd",x"8d",x"2c",x"d2",x"8a",x"1c",x"e7",
	x"fe",x"24",x"f5",x"20",x"01",x"e7",x"fe",x"28",x"20",x"12",x"e7",x"fe",x"29",x"28",x"10",x"cd",
	x"fb",x"24",x"df",x"fe",x"2c",x"20",x"03",x"e7",x"18",x"f5",x"fe",x"29",x"c2",x"8a",x"1c",x"e7",
	x"21",x"3b",x"5c",x"cb",x"b6",x"f1",x"28",x"02",x"cb",x"f6",x"c3",x"12",x"27",x"e7",x"e6",x"df",
	x"47",x"e7",x"d6",x"24",x"4f",x"20",x"01",x"e7",x"e7",x"e5",x"2a",x"53",x"5c",x"2b",x"11",x"ce",
	x"00",x"c5",x"cd",x"86",x"1d",x"c1",x"30",x"02",x"cf",x"18",x"e5",x"cd",x"ab",x"28",x"e6",x"df",
	x"b8",x"20",x"08",x"cd",x"ab",x"28",x"d6",x"24",x"b9",x"28",x"0c",x"e1",x"2b",x"11",x"00",x"02",
	x"c5",x"cd",x"8b",x"19",x"c1",x"18",x"d7",x"a7",x"cc",x"ab",x"28",x"d1",x"d1",x"ed",x"53",x"5d",
	x"5c",x"cd",x"ab",x"28",x"e5",x"fe",x"29",x"28",x"42",x"23",x"7e",x"fe",x"0e",x"16",x"40",x"28",
	x"07",x"2b",x"cd",x"ab",x"28",x"23",x"16",x"00",x"23",x"e5",x"d5",x"cd",x"fb",x"24",x"f1",x"fd",
	x"ae",x"01",x"e6",x"40",x"20",x"2b",x"e1",x"eb",x"2a",x"65",x"5c",x"01",x"05",x"00",x"ed",x"42",
	x"22",x"65",x"5c",x"ed",x"b0",x"eb",x"2b",x"cd",x"ab",x"28",x"fe",x"29",x"28",x"0d",x"e5",x"df",
	x"fe",x"2c",x"20",x"0d",x"e7",x"e1",x"cd",x"ab",x"28",x"18",x"be",x"e5",x"df",x"fe",x"29",x"28",
	x"02",x"cf",x"19",x"d1",x"eb",x"22",x"5d",x"5c",x"2a",x"0b",x"5c",x"e3",x"22",x"0b",x"5c",x"d5",
	x"e7",x"e7",x"cd",x"fb",x"24",x"e1",x"22",x"5d",x"5c",x"e1",x"22",x"0b",x"5c",x"e7",x"c3",x"12",
	x"27",x"23",x"7e",x"fe",x"21",x"38",x"fa",x"c9",x"fd",x"cb",x"01",x"f6",x"df",x"cd",x"8d",x"2c",
	x"d2",x"8a",x"1c",x"e5",x"e6",x"1f",x"4f",x"e7",x"e5",x"fe",x"28",x"28",x"28",x"cb",x"f1",x"fe",
	x"24",x"28",x"11",x"cb",x"e9",x"cd",x"88",x"2c",x"30",x"0f",x"cd",x"88",x"2c",x"30",x"16",x"cb",
	x"b1",x"e7",x"18",x"f6",x"e7",x"fd",x"cb",x"01",x"b6",x"3a",x"0c",x"5c",x"a7",x"28",x"06",x"cd",
	x"30",x"25",x"c2",x"51",x"29",x"41",x"cd",x"30",x"25",x"20",x"08",x"79",x"e6",x"e0",x"cb",x"ff",
	x"4f",x"18",x"37",x"2a",x"4b",x"5c",x"7e",x"e6",x"7f",x"28",x"2d",x"b9",x"20",x"22",x"17",x"87",
	x"f2",x"3f",x"29",x"38",x"30",x"d1",x"d5",x"e5",x"23",x"1a",x"13",x"fe",x"20",x"28",x"fa",x"f6",
	x"20",x"be",x"28",x"f4",x"f6",x"80",x"be",x"20",x"06",x"1a",x"cd",x"88",x"2c",x"30",x"15",x"e1",
	x"c5",x"cd",x"b8",x"19",x"eb",x"c1",x"18",x"ce",x"cb",x"f8",x"d1",x"df",x"fe",x"28",x"28",x"09",
	x"cb",x"e8",x"18",x"0d",x"d1",x"d1",x"d1",x"e5",x"df",x"cd",x"88",x"2c",x"30",x"03",x"e7",x"18",
	x"f8",x"e1",x"cb",x"10",x"cb",x"70",x"c9",x"2a",x"0b",x"5c",x"7e",x"fe",x"29",x"ca",x"ef",x"28",
	x"7e",x"f6",x"60",x"47",x"23",x"7e",x"fe",x"0e",x"28",x"07",x"2b",x"cd",x"ab",x"28",x"23",x"cb",
	x"a8",x"78",x"b9",x"28",x"12",x"23",x"23",x"23",x"23",x"23",x"cd",x"ab",x"28",x"fe",x"29",x"ca",
	x"ef",x"28",x"cd",x"ab",x"28",x"18",x"d9",x"cb",x"69",x"20",x"0c",x"23",x"ed",x"5b",x"65",x"5c",
	x"cd",x"c0",x"33",x"eb",x"22",x"65",x"5c",x"d1",x"d1",x"af",x"3c",x"c9",x"af",x"47",x"cb",x"79",
	x"20",x"4b",x"cb",x"7e",x"20",x"0e",x"3c",x"23",x"4e",x"23",x"46",x"23",x"eb",x"cd",x"b2",x"2a",
	x"df",x"c3",x"49",x"2a",x"23",x"23",x"23",x"46",x"cb",x"71",x"28",x"0a",x"05",x"28",x"e8",x"eb",
	x"df",x"fe",x"28",x"20",x"61",x"eb",x"eb",x"18",x"24",x"e5",x"df",x"e1",x"fe",x"2c",x"28",x"20",
	x"cb",x"79",x"28",x"52",x"cb",x"71",x"20",x"06",x"fe",x"29",x"20",x"3c",x"e7",x"c9",x"fe",x"29",
	x"28",x"6c",x"fe",x"cc",x"20",x"32",x"df",x"2b",x"22",x"5d",x"5c",x"18",x"5e",x"21",x"00",x"00",
	x"e5",x"e7",x"e1",x"79",x"fe",x"c0",x"20",x"09",x"df",x"fe",x"29",x"28",x"51",x"fe",x"cc",x"28",
	x"e5",x"c5",x"e5",x"cd",x"ee",x"2a",x"e3",x"eb",x"cd",x"cc",x"2a",x"38",x"19",x"0b",x"cd",x"f4",
	x"2a",x"09",x"d1",x"c1",x"10",x"b3",x"cb",x"79",x"20",x"66",x"e5",x"cb",x"71",x"20",x"13",x"42",
	x"4b",x"df",x"fe",x"29",x"28",x"02",x"cf",x"02",x"e7",x"e1",x"11",x"05",x"00",x"cd",x"f4",x"2a",
	x"09",x"c9",x"cd",x"ee",x"2a",x"e3",x"cd",x"f4",x"2a",x"c1",x"09",x"23",x"42",x"4b",x"eb",x"cd",
	x"b1",x"2a",x"df",x"fe",x"29",x"28",x"07",x"fe",x"2c",x"20",x"db",x"cd",x"52",x"2a",x"e7",x"fe",
	x"28",x"28",x"f8",x"fd",x"cb",x"01",x"b6",x"c9",x"cd",x"30",x"25",x"c4",x"f1",x"2b",x"e7",x"fe",
	x"29",x"28",x"50",x"d5",x"af",x"f5",x"c5",x"11",x"01",x"00",x"df",x"e1",x"fe",x"cc",x"28",x"17",
	x"f1",x"cd",x"cd",x"2a",x"f5",x"50",x"59",x"e5",x"df",x"e1",x"fe",x"cc",x"28",x"09",x"fe",x"29",
	x"c2",x"8a",x"1c",x"62",x"6b",x"18",x"13",x"e5",x"e7",x"e1",x"fe",x"29",x"28",x"0c",x"f1",x"cd",
	x"cd",x"2a",x"f5",x"df",x"60",x"69",x"fe",x"29",x"20",x"e6",x"f1",x"e3",x"19",x"2b",x"e3",x"a7",
	x"ed",x"52",x"01",x"00",x"00",x"38",x"07",x"23",x"a7",x"fa",x"20",x"2a",x"44",x"4d",x"d1",x"fd",
	x"cb",x"01",x"b6",x"cd",x"30",x"25",x"c8",x"af",x"fd",x"cb",x"01",x"b6",x"c5",x"cd",x"a9",x"33",
	x"c1",x"2a",x"65",x"5c",x"77",x"23",x"73",x"23",x"72",x"23",x"71",x"23",x"70",x"23",x"22",x"65",
	x"5c",x"c9",x"af",x"d5",x"e5",x"f5",x"cd",x"82",x"1c",x"f1",x"cd",x"30",x"25",x"28",x"12",x"f5",
	x"cd",x"99",x"1e",x"d1",x"78",x"b1",x"37",x"28",x"05",x"e1",x"e5",x"a7",x"ed",x"42",x"7a",x"de",
	x"00",x"e1",x"d1",x"c9",x"eb",x"23",x"5e",x"23",x"56",x"c9",x"cd",x"30",x"25",x"c8",x"cd",x"a9",
	x"30",x"da",x"15",x"1f",x"c9",x"2a",x"4d",x"5c",x"fd",x"cb",x"37",x"4e",x"28",x"5e",x"01",x"05",
	x"00",x"03",x"23",x"7e",x"fe",x"20",x"28",x"fa",x"30",x"0b",x"fe",x"10",x"38",x"11",x"fe",x"16",
	x"30",x"0d",x"23",x"18",x"ed",x"cd",x"88",x"2c",x"38",x"e7",x"fe",x"24",x"ca",x"c0",x"2b",x"79",
	x"2a",x"59",x"5c",x"2b",x"cd",x"55",x"16",x"23",x"23",x"eb",x"d5",x"2a",x"4d",x"5c",x"1b",x"d6",
	x"06",x"47",x"28",x"11",x"23",x"7e",x"fe",x"21",x"38",x"fa",x"f6",x"20",x"13",x"12",x"10",x"f4",
	x"f6",x"80",x"12",x"3e",x"c0",x"2a",x"4d",x"5c",x"ae",x"f6",x"20",x"e1",x"cd",x"ea",x"2b",x"e5",
	x"ef",x"02",x"38",x"e1",x"01",x"05",x"00",x"a7",x"ed",x"42",x"18",x"40",x"fd",x"cb",x"01",x"76",
	x"28",x"06",x"11",x"06",x"00",x"19",x"18",x"e7",x"2a",x"4d",x"5c",x"ed",x"4b",x"72",x"5c",x"fd",
	x"cb",x"37",x"46",x"20",x"30",x"78",x"b1",x"c8",x"e5",x"f7",x"d5",x"c5",x"54",x"5d",x"23",x"36",
	x"20",x"ed",x"b8",x"e5",x"cd",x"f1",x"2b",x"e1",x"e3",x"a7",x"ed",x"42",x"09",x"30",x"02",x"44",
	x"4d",x"e3",x"eb",x"78",x"b1",x"28",x"02",x"ed",x"b0",x"c1",x"d1",x"e1",x"eb",x"78",x"b1",x"c8",
	x"d5",x"ed",x"b0",x"e1",x"c9",x"2b",x"2b",x"2b",x"7e",x"e5",x"c5",x"cd",x"c6",x"2b",x"c1",x"e1",
	x"03",x"03",x"03",x"c3",x"e8",x"19",x"3e",x"df",x"2a",x"4d",x"5c",x"a6",x"f5",x"cd",x"f1",x"2b",
	x"eb",x"09",x"c5",x"2b",x"22",x"4d",x"5c",x"03",x"03",x"03",x"2a",x"59",x"5c",x"2b",x"cd",x"55",
	x"16",x"2a",x"4d",x"5c",x"c1",x"c5",x"03",x"ed",x"b8",x"eb",x"23",x"c1",x"70",x"2b",x"71",x"f1",
	x"2b",x"77",x"2a",x"59",x"5c",x"2b",x"c9",x"2a",x"65",x"5c",x"2b",x"46",x"2b",x"4e",x"2b",x"56",
	x"2b",x"5e",x"2b",x"7e",x"22",x"65",x"5c",x"c9",x"cd",x"b2",x"28",x"c2",x"8a",x"1c",x"cd",x"30",
	x"25",x"20",x"08",x"cb",x"b1",x"cd",x"96",x"29",x"cd",x"ee",x"1b",x"38",x"08",x"c5",x"cd",x"b8",
	x"19",x"cd",x"e8",x"19",x"c1",x"cb",x"f9",x"06",x"00",x"c5",x"21",x"01",x"00",x"cb",x"71",x"20",
	x"02",x"2e",x"05",x"eb",x"e7",x"26",x"ff",x"cd",x"cc",x"2a",x"da",x"20",x"2a",x"e1",x"c5",x"24",
	x"e5",x"60",x"69",x"cd",x"f4",x"2a",x"eb",x"df",x"fe",x"2c",x"28",x"e8",x"fe",x"29",x"20",x"bb",
	x"e7",x"c1",x"79",x"68",x"26",x"00",x"23",x"23",x"29",x"19",x"da",x"15",x"1f",x"d5",x"c5",x"e5",
	x"44",x"4d",x"2a",x"59",x"5c",x"2b",x"cd",x"55",x"16",x"23",x"77",x"c1",x"0b",x"0b",x"0b",x"23",
	x"71",x"23",x"70",x"c1",x"78",x"23",x"77",x"62",x"6b",x"1b",x"36",x"00",x"cb",x"71",x"28",x"02",
	x"36",x"20",x"c1",x"ed",x"b8",x"c1",x"70",x"2b",x"71",x"2b",x"3d",x"20",x"f8",x"c9",x"cd",x"1b",
	x"2d",x"3f",x"d8",x"fe",x"41",x"3f",x"d0",x"fe",x"5b",x"d8",x"fe",x"61",x"3f",x"d0",x"fe",x"7b",
	x"c9",x"fe",x"c4",x"20",x"19",x"11",x"00",x"00",x"e7",x"d6",x"31",x"ce",x"00",x"20",x"0a",x"eb",
	x"3f",x"ed",x"6a",x"da",x"ad",x"31",x"eb",x"18",x"ef",x"42",x"4b",x"c3",x"2b",x"2d",x"fe",x"2e",
	x"28",x"0f",x"cd",x"3b",x"2d",x"fe",x"2e",x"20",x"28",x"e7",x"cd",x"1b",x"2d",x"38",x"22",x"18",
	x"0a",x"e7",x"cd",x"1b",x"2d",x"da",x"8a",x"1c",x"ef",x"a0",x"38",x"ef",x"a1",x"c0",x"02",x"38",
	x"df",x"cd",x"22",x"2d",x"38",x"0b",x"ef",x"e0",x"a4",x"05",x"c0",x"04",x"0f",x"38",x"e7",x"18",
	x"ef",x"fe",x"45",x"28",x"03",x"fe",x"65",x"c0",x"06",x"ff",x"e7",x"fe",x"2b",x"28",x"05",x"fe",
	x"2d",x"20",x"02",x"04",x"e7",x"cd",x"1b",x"2d",x"38",x"cb",x"c5",x"cd",x"3b",x"2d",x"cd",x"d5",
	x"2d",x"c1",x"da",x"ad",x"31",x"a7",x"fa",x"ad",x"31",x"04",x"28",x"02",x"ed",x"44",x"c3",x"4f",
	x"2d",x"fe",x"30",x"d8",x"fe",x"3a",x"3f",x"c9",x"cd",x"1b",x"2d",x"d8",x"d6",x"30",x"4f",x"06",
	x"00",x"fd",x"21",x"3a",x"5c",x"af",x"5f",x"51",x"48",x"47",x"cd",x"b6",x"2a",x"ef",x"38",x"a7",
	x"c9",x"f5",x"ef",x"a0",x"38",x"f1",x"cd",x"22",x"2d",x"d8",x"ef",x"01",x"a4",x"04",x"0f",x"38",
	x"cd",x"74",x"00",x"18",x"f1",x"07",x"0f",x"30",x"02",x"2f",x"3c",x"f5",x"21",x"92",x"5c",x"cd",
	x"0b",x"35",x"ef",x"a4",x"38",x"f1",x"cb",x"3f",x"30",x"0d",x"f5",x"ef",x"c1",x"e0",x"00",x"04",
	x"04",x"33",x"02",x"05",x"e1",x"38",x"f1",x"28",x"08",x"f5",x"ef",x"31",x"04",x"38",x"f1",x"18",
	x"e5",x"ef",x"02",x"38",x"c9",x"23",x"4e",x"23",x"7e",x"a9",x"91",x"5f",x"23",x"7e",x"89",x"a9",
	x"57",x"c9",x"0e",x"00",x"e5",x"36",x"00",x"23",x"71",x"23",x"7b",x"a9",x"91",x"77",x"23",x"7a",
	x"89",x"a9",x"77",x"23",x"36",x"00",x"e1",x"c9",x"ef",x"38",x"7e",x"a7",x"28",x"05",x"ef",x"a2",
	x"0f",x"27",x"38",x"ef",x"02",x"38",x"e5",x"d5",x"eb",x"46",x"cd",x"7f",x"2d",x"af",x"90",x"cb",
	x"79",x"42",x"4b",x"7b",x"d1",x"e1",x"c9",x"57",x"17",x"9f",x"5f",x"4f",x"af",x"47",x"cd",x"b6",
	x"2a",x"ef",x"34",x"ef",x"1a",x"20",x"9a",x"85",x"04",x"27",x"38",x"cd",x"a2",x"2d",x"d8",x"f5",
	x"05",x"04",x"28",x"03",x"f1",x"37",x"c9",x"f1",x"c9",x"ef",x"31",x"36",x"00",x"0b",x"31",x"37",
	x"00",x"0d",x"02",x"38",x"3e",x"30",x"d7",x"c9",x"2a",x"38",x"3e",x"2d",x"d7",x"ef",x"a0",x"c3",
	x"c4",x"c5",x"02",x"38",x"d9",x"e5",x"d9",x"ef",x"31",x"27",x"c2",x"03",x"e2",x"01",x"c2",x"02",
	x"38",x"7e",x"a7",x"20",x"47",x"cd",x"7f",x"2d",x"06",x"10",x"7a",x"a7",x"20",x"06",x"b3",x"28",
	x"09",x"53",x"06",x"08",x"d5",x"d9",x"d1",x"d9",x"18",x"57",x"ef",x"e2",x"38",x"7e",x"d6",x"7e",
	x"cd",x"c1",x"2d",x"57",x"3a",x"ac",x"5c",x"92",x"32",x"ac",x"5c",x"7a",x"cd",x"4f",x"2d",x"ef",
	x"31",x"27",x"c1",x"03",x"e1",x"38",x"cd",x"d5",x"2d",x"e5",x"32",x"a1",x"5c",x"3d",x"17",x"9f",
	x"3c",x"21",x"ab",x"5c",x"77",x"23",x"86",x"77",x"e1",x"c3",x"cf",x"2e",x"d6",x"80",x"fe",x"1c",
	x"38",x"13",x"cd",x"c1",x"2d",x"d6",x"07",x"47",x"21",x"ac",x"5c",x"86",x"77",x"78",x"ed",x"44",
	x"cd",x"4f",x"2d",x"18",x"92",x"eb",x"cd",x"ba",x"2f",x"d9",x"cb",x"fa",x"7d",x"d9",x"d6",x"80",
	x"47",x"cb",x"23",x"cb",x"12",x"d9",x"cb",x"13",x"cb",x"12",x"d9",x"21",x"aa",x"5c",x"0e",x"05",
	x"7e",x"8f",x"27",x"77",x"2b",x"0d",x"20",x"f8",x"10",x"e7",x"af",x"21",x"a6",x"5c",x"11",x"a1",
	x"5c",x"06",x"09",x"ed",x"6f",x"0e",x"ff",x"ed",x"6f",x"20",x"04",x"0d",x"0c",x"20",x"0a",x"12",
	x"13",x"fd",x"34",x"71",x"fd",x"34",x"72",x"0e",x"00",x"cb",x"40",x"28",x"01",x"23",x"10",x"e7",
	x"3a",x"ab",x"5c",x"d6",x"09",x"38",x"0a",x"fd",x"35",x"71",x"3e",x"04",x"fd",x"be",x"6f",x"18",
	x"41",x"ef",x"02",x"e2",x"38",x"eb",x"cd",x"ba",x"2f",x"d9",x"3e",x"80",x"95",x"2e",x"00",x"cb",
	x"fa",x"d9",x"cd",x"dd",x"2f",x"fd",x"7e",x"71",x"fe",x"08",x"38",x"06",x"d9",x"cb",x"12",x"d9",
	x"18",x"20",x"01",x"00",x"02",x"7b",x"cd",x"8b",x"2f",x"5f",x"7a",x"cd",x"8b",x"2f",x"57",x"c5",
	x"d9",x"c1",x"10",x"f1",x"21",x"a1",x"5c",x"79",x"fd",x"4e",x"71",x"09",x"77",x"fd",x"34",x"71",
	x"18",x"d3",x"f5",x"21",x"a1",x"5c",x"fd",x"4e",x"71",x"06",x"00",x"09",x"41",x"f1",x"2b",x"7e",
	x"ce",x"00",x"77",x"a7",x"28",x"05",x"fe",x"0a",x"3f",x"30",x"08",x"10",x"f1",x"36",x"01",x"04",
	x"fd",x"34",x"72",x"fd",x"70",x"71",x"ef",x"02",x"38",x"d9",x"e1",x"d9",x"ed",x"4b",x"ab",x"5c",
	x"21",x"a1",x"5c",x"78",x"fe",x"09",x"38",x"04",x"fe",x"fc",x"38",x"26",x"a7",x"cc",x"ef",x"15",
	x"af",x"90",x"fa",x"52",x"2f",x"47",x"18",x"0c",x"79",x"a7",x"28",x"03",x"7e",x"23",x"0d",x"cd",
	x"ef",x"15",x"10",x"f4",x"79",x"a7",x"c8",x"04",x"3e",x"2e",x"d7",x"3e",x"30",x"10",x"fb",x"41",
	x"18",x"e6",x"50",x"15",x"06",x"01",x"cd",x"4a",x"2f",x"3e",x"45",x"d7",x"4a",x"79",x"a7",x"f2",
	x"83",x"2f",x"ed",x"44",x"4f",x"3e",x"2d",x"18",x"02",x"3e",x"2b",x"d7",x"06",x"00",x"c3",x"1b",
	x"1a",x"d5",x"6f",x"26",x"00",x"5d",x"54",x"29",x"29",x"19",x"29",x"59",x"19",x"4c",x"7d",x"d1",
	x"c9",x"7e",x"36",x"00",x"a7",x"c8",x"23",x"cb",x"7e",x"cb",x"fe",x"2b",x"c8",x"c5",x"01",x"05",
	x"00",x"09",x"41",x"4f",x"37",x"2b",x"7e",x"2f",x"ce",x"00",x"77",x"10",x"f8",x"79",x"c1",x"c9",
	x"e5",x"f5",x"4e",x"23",x"46",x"77",x"23",x"79",x"4e",x"c5",x"23",x"4e",x"23",x"46",x"eb",x"57",
	x"5e",x"d5",x"23",x"56",x"23",x"5e",x"d5",x"d9",x"d1",x"e1",x"c1",x"d9",x"23",x"56",x"23",x"5e",
	x"f1",x"e1",x"c9",x"a7",x"c8",x"fe",x"21",x"30",x"16",x"c5",x"47",x"d9",x"cb",x"2d",x"cb",x"1a",
	x"cb",x"1b",x"d9",x"cb",x"1a",x"cb",x"1b",x"10",x"f2",x"c1",x"d0",x"cd",x"04",x"30",x"c0",x"d9",
	x"af",x"2e",x"00",x"57",x"5d",x"d9",x"11",x"00",x"00",x"c9",x"1c",x"c0",x"14",x"c0",x"d9",x"1c",
	x"20",x"01",x"14",x"d9",x"c9",x"eb",x"cd",x"6e",x"34",x"eb",x"1a",x"b6",x"20",x"26",x"d5",x"23",
	x"e5",x"23",x"5e",x"23",x"56",x"23",x"23",x"23",x"7e",x"23",x"4e",x"23",x"46",x"e1",x"eb",x"09",
	x"eb",x"8e",x"0f",x"ce",x"00",x"20",x"0b",x"9f",x"77",x"23",x"73",x"23",x"72",x"2b",x"2b",x"2b",
	x"d1",x"c9",x"2b",x"d1",x"cd",x"93",x"32",x"d9",x"e5",x"d9",x"d5",x"e5",x"cd",x"9b",x"2f",x"47",
	x"eb",x"cd",x"9b",x"2f",x"4f",x"b8",x"30",x"03",x"78",x"41",x"eb",x"f5",x"90",x"cd",x"ba",x"2f",
	x"cd",x"dd",x"2f",x"f1",x"e1",x"77",x"e5",x"68",x"61",x"19",x"d9",x"eb",x"ed",x"4a",x"eb",x"7c",
	x"8d",x"6f",x"1f",x"ad",x"d9",x"eb",x"e1",x"1f",x"30",x"08",x"3e",x"01",x"cd",x"dd",x"2f",x"34",
	x"28",x"23",x"d9",x"7d",x"e6",x"80",x"d9",x"23",x"77",x"2b",x"28",x"1f",x"7b",x"ed",x"44",x"3f",
	x"5f",x"7a",x"2f",x"ce",x"00",x"57",x"d9",x"7b",x"2f",x"ce",x"00",x"5f",x"7a",x"2f",x"ce",x"00",
	x"30",x"07",x"1f",x"d9",x"34",x"ca",x"ad",x"31",x"d9",x"57",x"d9",x"af",x"c3",x"55",x"31",x"c5",
	x"06",x"10",x"7c",x"4d",x"21",x"00",x"00",x"29",x"38",x"0a",x"cb",x"11",x"17",x"30",x"03",x"19",
	x"38",x"02",x"10",x"f3",x"c1",x"c9",x"cd",x"e9",x"34",x"d8",x"23",x"ae",x"cb",x"fe",x"2b",x"c9",
	x"1a",x"b6",x"20",x"22",x"d5",x"e5",x"d5",x"cd",x"7f",x"2d",x"eb",x"e3",x"41",x"cd",x"7f",x"2d",
	x"78",x"a9",x"4f",x"e1",x"cd",x"a9",x"30",x"eb",x"e1",x"38",x"0a",x"7a",x"b3",x"20",x"01",x"4f",
	x"cd",x"8e",x"2d",x"d1",x"c9",x"d1",x"cd",x"93",x"32",x"af",x"cd",x"c0",x"30",x"d8",x"d9",x"e5",
	x"d9",x"d5",x"eb",x"cd",x"c0",x"30",x"eb",x"38",x"5a",x"e5",x"cd",x"ba",x"2f",x"78",x"a7",x"ed",
	x"62",x"d9",x"e5",x"ed",x"62",x"d9",x"06",x"21",x"18",x"11",x"30",x"05",x"19",x"d9",x"ed",x"5a",
	x"d9",x"d9",x"cb",x"1c",x"cb",x"1d",x"d9",x"cb",x"1c",x"cb",x"1d",x"d9",x"cb",x"18",x"cb",x"19",
	x"d9",x"cb",x"19",x"1f",x"10",x"e4",x"eb",x"d9",x"eb",x"d9",x"c1",x"e1",x"78",x"81",x"20",x"01",
	x"a7",x"3d",x"3f",x"17",x"3f",x"1f",x"f2",x"46",x"31",x"30",x"68",x"a7",x"3c",x"20",x"08",x"38",
	x"06",x"d9",x"cb",x"7a",x"d9",x"20",x"5c",x"77",x"d9",x"78",x"d9",x"30",x"15",x"7e",x"a7",x"3e",
	x"80",x"28",x"01",x"af",x"d9",x"a2",x"cd",x"fb",x"2f",x"07",x"77",x"38",x"2e",x"23",x"77",x"2b",
	x"18",x"29",x"06",x"20",x"d9",x"cb",x"7a",x"d9",x"20",x"12",x"07",x"cb",x"13",x"cb",x"12",x"d9",
	x"cb",x"13",x"cb",x"12",x"d9",x"35",x"28",x"d7",x"10",x"ea",x"18",x"d7",x"17",x"30",x"0c",x"cd",
	x"04",x"30",x"20",x"07",x"d9",x"16",x"80",x"d9",x"34",x"28",x"18",x"e5",x"23",x"d9",x"d5",x"d9",
	x"c1",x"78",x"17",x"cb",x"16",x"1f",x"77",x"23",x"71",x"23",x"72",x"23",x"73",x"e1",x"d1",x"d9",
	x"e1",x"d9",x"c9",x"cf",x"05",x"cd",x"93",x"32",x"eb",x"af",x"cd",x"c0",x"30",x"38",x"f4",x"eb",
	x"cd",x"c0",x"30",x"d8",x"d9",x"e5",x"d9",x"d5",x"e5",x"cd",x"ba",x"2f",x"d9",x"e5",x"60",x"69",
	x"d9",x"61",x"68",x"af",x"06",x"df",x"18",x"10",x"17",x"cb",x"11",x"d9",x"cb",x"11",x"cb",x"10",
	x"d9",x"29",x"d9",x"ed",x"6a",x"d9",x"38",x"10",x"ed",x"52",x"d9",x"ed",x"52",x"d9",x"30",x"0f",
	x"19",x"d9",x"ed",x"5a",x"d9",x"a7",x"18",x"08",x"a7",x"ed",x"52",x"d9",x"ed",x"52",x"d9",x"37",
	x"04",x"fa",x"d2",x"31",x"f5",x"28",x"e1",x"5f",x"51",x"d9",x"59",x"50",x"f1",x"cb",x"18",x"f1",
	x"cb",x"18",x"d9",x"c1",x"e1",x"78",x"91",x"c3",x"3d",x"31",x"7e",x"a7",x"c8",x"fe",x"81",x"30",
	x"06",x"36",x"00",x"3e",x"20",x"18",x"51",x"fe",x"91",x"20",x"1a",x"23",x"23",x"23",x"3e",x"80",
	x"a6",x"2b",x"b6",x"2b",x"20",x"03",x"3e",x"80",x"ae",x"2b",x"20",x"36",x"77",x"23",x"36",x"ff",
	x"2b",x"3e",x"18",x"18",x"33",x"30",x"2c",x"d5",x"2f",x"c6",x"91",x"23",x"56",x"23",x"5e",x"2b",
	x"2b",x"0e",x"00",x"cb",x"7a",x"28",x"01",x"0d",x"cb",x"fa",x"06",x"08",x"90",x"80",x"38",x"04",
	x"5a",x"16",x"00",x"90",x"28",x"07",x"47",x"cb",x"3a",x"cb",x"1b",x"10",x"fa",x"cd",x"8e",x"2d",
	x"d1",x"c9",x"7e",x"d6",x"a0",x"f0",x"ed",x"44",x"d5",x"eb",x"2b",x"47",x"cb",x"38",x"cb",x"38",
	x"cb",x"38",x"28",x"05",x"36",x"00",x"2b",x"10",x"fb",x"e6",x"07",x"28",x"09",x"47",x"3e",x"ff",
	x"cb",x"27",x"10",x"fc",x"a6",x"77",x"eb",x"d1",x"c9",x"cd",x"96",x"32",x"eb",x"7e",x"a7",x"c0",
	x"d5",x"cd",x"7f",x"2d",x"af",x"23",x"77",x"2b",x"77",x"06",x"91",x"7a",x"a7",x"20",x"08",x"b3",
	x"42",x"28",x"10",x"53",x"58",x"06",x"89",x"eb",x"05",x"29",x"30",x"fc",x"cb",x"09",x"cb",x"1c",
	x"cb",x"1d",x"eb",x"2b",x"73",x"2b",x"72",x"2b",x"70",x"d1",x"c9",x"00",x"b0",x"00",x"40",x"b0",
	x"00",x"01",x"30",x"00",x"f1",x"49",x"0f",x"da",x"a2",x"40",x"b0",x"00",x"0a",x"8f",x"36",x"3c",
	x"34",x"a1",x"33",x"0f",x"30",x"ca",x"30",x"af",x"31",x"51",x"38",x"1b",x"35",x"24",x"35",x"3b",
	x"35",x"3b",x"35",x"3b",x"35",x"3b",x"35",x"3b",x"35",x"3b",x"35",x"14",x"30",x"2d",x"35",x"3b",
	x"35",x"3b",x"35",x"3b",x"35",x"3b",x"35",x"3b",x"35",x"3b",x"35",x"9c",x"35",x"de",x"35",x"bc",
	x"34",x"45",x"36",x"6e",x"34",x"69",x"36",x"de",x"35",x"74",x"36",x"b5",x"37",x"aa",x"37",x"da",
	x"37",x"33",x"38",x"43",x"38",x"e2",x"37",x"13",x"37",x"c4",x"36",x"af",x"36",x"4a",x"38",x"92",
	x"34",x"6a",x"34",x"ac",x"34",x"a5",x"34",x"b3",x"34",x"1f",x"36",x"c9",x"35",x"01",x"35",x"c0",
	x"33",x"a0",x"36",x"86",x"36",x"c6",x"33",x"7a",x"36",x"06",x"35",x"f9",x"34",x"9b",x"36",x"83",
	x"37",x"14",x"32",x"a2",x"33",x"4f",x"2d",x"97",x"32",x"49",x"34",x"1b",x"34",x"2d",x"34",x"0f",
	x"34",x"cd",x"bf",x"35",x"78",x"32",x"67",x"5c",x"d9",x"e3",x"d9",x"ed",x"53",x"65",x"5c",x"d9",
	x"7e",x"23",x"e5",x"a7",x"f2",x"80",x"33",x"57",x"e6",x"60",x"0f",x"0f",x"0f",x"0f",x"c6",x"7c",
	x"6f",x"7a",x"e6",x"1f",x"18",x"0e",x"fe",x"18",x"30",x"08",x"d9",x"01",x"fb",x"ff",x"54",x"5d",
	x"09",x"d9",x"07",x"6f",x"11",x"d7",x"32",x"26",x"00",x"19",x"5e",x"23",x"56",x"21",x"65",x"33",
	x"e3",x"d5",x"d9",x"ed",x"4b",x"66",x"5c",x"c9",x"f1",x"3a",x"67",x"5c",x"d9",x"18",x"c3",x"d5",
	x"e5",x"01",x"05",x"00",x"cd",x"05",x"1f",x"e1",x"d1",x"c9",x"ed",x"5b",x"65",x"5c",x"cd",x"c0",
	x"33",x"ed",x"53",x"65",x"5c",x"c9",x"cd",x"a9",x"33",x"ed",x"b0",x"c9",x"62",x"6b",x"cd",x"a9",
	x"33",x"d9",x"e5",x"d9",x"e3",x"c5",x"7e",x"e6",x"c0",x"07",x"07",x"4f",x"0c",x"7e",x"e6",x"3f",
	x"20",x"02",x"23",x"7e",x"c6",x"50",x"12",x"3e",x"05",x"91",x"23",x"13",x"06",x"00",x"ed",x"b0",
	x"c1",x"e3",x"d9",x"e1",x"d9",x"47",x"af",x"05",x"c8",x"12",x"13",x"18",x"fa",x"a7",x"c8",x"f5",
	x"d5",x"11",x"00",x"00",x"cd",x"c8",x"33",x"d1",x"f1",x"3d",x"18",x"f2",x"4f",x"07",x"07",x"81",
	x"4f",x"06",x"00",x"09",x"c9",x"d5",x"2a",x"68",x"5c",x"cd",x"06",x"34",x"cd",x"c0",x"33",x"e1",
	x"c9",x"62",x"6b",x"d9",x"e5",x"21",x"c5",x"32",x"d9",x"cd",x"f7",x"33",x"cd",x"c8",x"33",x"d9",
	x"e1",x"d9",x"c9",x"e5",x"eb",x"2a",x"68",x"5c",x"cd",x"06",x"34",x"eb",x"cd",x"c0",x"33",x"eb",
	x"e1",x"c9",x"06",x"05",x"1a",x"4e",x"eb",x"12",x"71",x"23",x"13",x"10",x"f7",x"eb",x"c9",x"47",
	x"cd",x"5e",x"33",x"31",x"0f",x"c0",x"02",x"a0",x"c2",x"31",x"e0",x"04",x"e2",x"c1",x"03",x"38",
	x"cd",x"c6",x"33",x"cd",x"62",x"33",x"0f",x"01",x"c2",x"02",x"35",x"ee",x"e1",x"03",x"38",x"c9",
	x"06",x"ff",x"18",x"06",x"cd",x"e9",x"34",x"d8",x"06",x"00",x"7e",x"a7",x"28",x"0b",x"23",x"78",
	x"e6",x"80",x"b6",x"17",x"3f",x"1f",x"77",x"2b",x"c9",x"d5",x"e5",x"cd",x"7f",x"2d",x"e1",x"78",
	x"b1",x"2f",x"4f",x"cd",x"8e",x"2d",x"d1",x"c9",x"cd",x"e9",x"34",x"d8",x"d5",x"11",x"01",x"00",
	x"23",x"cb",x"16",x"2b",x"9f",x"4f",x"cd",x"8e",x"2d",x"d1",x"c9",x"cd",x"99",x"1e",x"ed",x"78",
	x"18",x"04",x"cd",x"99",x"1e",x"0a",x"c3",x"28",x"2d",x"cd",x"99",x"1e",x"21",x"2b",x"2d",x"e5",
	x"c5",x"c9",x"cd",x"f1",x"2b",x"0b",x"78",x"b1",x"20",x"23",x"1a",x"cd",x"8d",x"2c",x"38",x"09",
	x"d6",x"90",x"38",x"19",x"fe",x"15",x"30",x"15",x"3c",x"3d",x"87",x"87",x"87",x"fe",x"a8",x"30",
	x"0c",x"ed",x"4b",x"7b",x"5c",x"81",x"4f",x"30",x"01",x"04",x"c3",x"2b",x"2d",x"cf",x"09",x"e5",
	x"c5",x"47",x"7e",x"23",x"b6",x"23",x"b6",x"23",x"b6",x"78",x"c1",x"e1",x"c0",x"37",x"c9",x"cd",
	x"e9",x"34",x"d8",x"3e",x"ff",x"18",x"06",x"cd",x"e9",x"34",x"18",x"05",x"af",x"23",x"ae",x"2b",
	x"07",x"e5",x"3e",x"00",x"77",x"23",x"77",x"23",x"17",x"77",x"1f",x"23",x"77",x"23",x"77",x"e1",
	x"c9",x"eb",x"cd",x"e9",x"34",x"eb",x"d8",x"37",x"18",x"e7",x"eb",x"cd",x"e9",x"34",x"eb",x"d0",
	x"a7",x"18",x"de",x"eb",x"cd",x"e9",x"34",x"eb",x"d0",x"d5",x"1b",x"af",x"12",x"1b",x"12",x"d1",
	x"c9",x"78",x"d6",x"08",x"cb",x"57",x"20",x"01",x"3d",x"0f",x"30",x"08",x"f5",x"e5",x"cd",x"3c",
	x"34",x"d1",x"eb",x"f1",x"cb",x"57",x"20",x"07",x"0f",x"f5",x"cd",x"0f",x"30",x"18",x"33",x"0f",
	x"f5",x"cd",x"f1",x"2b",x"d5",x"c5",x"cd",x"f1",x"2b",x"e1",x"7c",x"b5",x"e3",x"78",x"20",x"0b",
	x"b1",x"c1",x"28",x"04",x"f1",x"3f",x"18",x"16",x"f1",x"18",x"13",x"b1",x"28",x"0d",x"1a",x"96",
	x"38",x"09",x"20",x"ed",x"0b",x"13",x"23",x"e3",x"2b",x"18",x"df",x"c1",x"f1",x"a7",x"f5",x"ef",
	x"a0",x"38",x"f1",x"f5",x"dc",x"01",x"35",x"f1",x"f5",x"d4",x"f9",x"34",x"f1",x"0f",x"d4",x"01",
	x"35",x"c9",x"cd",x"f1",x"2b",x"d5",x"c5",x"cd",x"f1",x"2b",x"e1",x"e5",x"d5",x"c5",x"09",x"44",
	x"4d",x"f7",x"cd",x"b2",x"2a",x"c1",x"e1",x"78",x"b1",x"28",x"02",x"ed",x"b0",x"c1",x"e1",x"78",
	x"b1",x"28",x"02",x"ed",x"b0",x"2a",x"65",x"5c",x"11",x"fb",x"ff",x"e5",x"19",x"d1",x"c9",x"cd",
	x"d5",x"2d",x"38",x"0e",x"20",x"0c",x"f5",x"01",x"01",x"00",x"f7",x"f1",x"12",x"cd",x"b2",x"2a",
	x"eb",x"c9",x"cf",x"0a",x"2a",x"5d",x"5c",x"e5",x"78",x"c6",x"e3",x"9f",x"f5",x"cd",x"f1",x"2b",
	x"d5",x"03",x"f7",x"e1",x"ed",x"53",x"5d",x"5c",x"d5",x"ed",x"b0",x"eb",x"2b",x"36",x"0d",x"fd",
	x"cb",x"01",x"be",x"cd",x"fb",x"24",x"df",x"fe",x"0d",x"20",x"07",x"e1",x"f1",x"fd",x"ae",x"01",
	x"e6",x"40",x"c2",x"8a",x"1c",x"22",x"5d",x"5c",x"fd",x"cb",x"01",x"fe",x"cd",x"fb",x"24",x"e1",
	x"22",x"5d",x"5c",x"18",x"a0",x"01",x"01",x"00",x"f7",x"22",x"5b",x"5c",x"e5",x"2a",x"51",x"5c",
	x"e5",x"3e",x"ff",x"cd",x"01",x"16",x"cd",x"e3",x"2d",x"e1",x"cd",x"15",x"16",x"d1",x"2a",x"5b",
	x"5c",x"a7",x"ed",x"52",x"44",x"4d",x"cd",x"b2",x"2a",x"eb",x"c9",x"cd",x"94",x"1e",x"fe",x"10",
	x"d2",x"9f",x"1e",x"2a",x"51",x"5c",x"e5",x"cd",x"01",x"16",x"cd",x"e6",x"15",x"01",x"00",x"00",
	x"30",x"03",x"0c",x"f7",x"12",x"cd",x"b2",x"2a",x"e1",x"cd",x"15",x"16",x"c3",x"bf",x"35",x"cd",
	x"f1",x"2b",x"78",x"b1",x"28",x"01",x"1a",x"c3",x"28",x"2d",x"cd",x"f1",x"2b",x"c3",x"2b",x"2d",
	x"d9",x"e5",x"21",x"67",x"5c",x"35",x"e1",x"20",x"04",x"23",x"d9",x"c9",x"d9",x"5e",x"7b",x"17",
	x"9f",x"57",x"19",x"d9",x"c9",x"13",x"13",x"1a",x"1b",x"1b",x"a7",x"20",x"ef",x"d9",x"23",x"d9",
	x"c9",x"f1",x"d9",x"e3",x"d9",x"c9",x"ef",x"c0",x"02",x"31",x"e0",x"05",x"27",x"e0",x"01",x"c0",
	x"04",x"03",x"e0",x"38",x"c9",x"ef",x"31",x"36",x"00",x"04",x"3a",x"38",x"c9",x"31",x"3a",x"c0",
	x"03",x"e0",x"01",x"30",x"00",x"03",x"a1",x"03",x"38",x"c9",x"ef",x"3d",x"34",x"f1",x"38",x"aa",
	x"3b",x"29",x"04",x"31",x"27",x"c3",x"03",x"31",x"0f",x"a1",x"03",x"88",x"13",x"36",x"58",x"65",
	x"66",x"9d",x"78",x"65",x"40",x"a2",x"60",x"32",x"c9",x"e7",x"21",x"f7",x"af",x"24",x"eb",x"2f",
	x"b0",x"b0",x"14",x"ee",x"7e",x"bb",x"94",x"58",x"f1",x"3a",x"7e",x"f8",x"cf",x"e3",x"38",x"cd",
	x"d5",x"2d",x"20",x"07",x"38",x"03",x"86",x"30",x"09",x"cf",x"05",x"38",x"07",x"96",x"30",x"04",
	x"ed",x"44",x"77",x"c9",x"ef",x"02",x"a0",x"38",x"c9",x"ef",x"3d",x"31",x"37",x"00",x"04",x"38",
	x"cf",x"09",x"a0",x"02",x"38",x"7e",x"36",x"80",x"cd",x"28",x"2d",x"ef",x"34",x"38",x"00",x"03",
	x"01",x"31",x"34",x"f0",x"4c",x"cc",x"cc",x"cd",x"03",x"37",x"00",x"08",x"01",x"a1",x"03",x"01",
	x"38",x"34",x"ef",x"01",x"34",x"f0",x"31",x"72",x"17",x"f8",x"04",x"01",x"a2",x"03",x"a2",x"03",
	x"31",x"34",x"32",x"20",x"04",x"a2",x"03",x"8c",x"11",x"ac",x"14",x"09",x"56",x"da",x"a5",x"59",
	x"30",x"c5",x"5c",x"90",x"aa",x"9e",x"70",x"6f",x"61",x"a1",x"cb",x"da",x"96",x"a4",x"31",x"9f",
	x"b4",x"e7",x"a0",x"fe",x"5c",x"fc",x"ea",x"1b",x"43",x"ca",x"36",x"ed",x"a7",x"9c",x"7e",x"5e",
	x"f0",x"6e",x"23",x"80",x"93",x"04",x"0f",x"38",x"c9",x"ef",x"3d",x"34",x"ee",x"22",x"f9",x"83",
	x"6e",x"04",x"31",x"a2",x"0f",x"27",x"03",x"31",x"0f",x"31",x"0f",x"31",x"2a",x"a1",x"03",x"31",
	x"37",x"c0",x"00",x"04",x"02",x"38",x"c9",x"a1",x"03",x"01",x"36",x"00",x"02",x"1b",x"38",x"c9",
	x"ef",x"39",x"2a",x"a1",x"03",x"e0",x"00",x"06",x"1b",x"33",x"03",x"ef",x"39",x"31",x"31",x"04",
	x"31",x"0f",x"a1",x"03",x"86",x"14",x"e6",x"5c",x"1f",x"0b",x"a3",x"8f",x"38",x"ee",x"e9",x"15",
	x"63",x"bb",x"23",x"ee",x"92",x"0d",x"cd",x"ed",x"f1",x"23",x"5d",x"1b",x"ea",x"04",x"38",x"c9",
	x"ef",x"31",x"1f",x"01",x"20",x"05",x"38",x"c9",x"cd",x"97",x"32",x"7e",x"fe",x"81",x"38",x"0e",
	x"ef",x"a1",x"1b",x"01",x"05",x"31",x"36",x"a3",x"01",x"00",x"06",x"1b",x"33",x"03",x"ef",x"a0",
	x"01",x"31",x"31",x"04",x"31",x"0f",x"a1",x"03",x"8c",x"10",x"b2",x"13",x"0e",x"55",x"e4",x"8d",
	x"58",x"39",x"bc",x"5b",x"98",x"fd",x"9e",x"00",x"36",x"75",x"a0",x"db",x"e8",x"b4",x"63",x"42",
	x"c4",x"e6",x"b5",x"09",x"36",x"be",x"e9",x"36",x"73",x"1b",x"5d",x"ec",x"d8",x"de",x"63",x"be",
	x"f0",x"61",x"a1",x"b3",x"0c",x"04",x"0f",x"38",x"c9",x"ef",x"31",x"31",x"04",x"a1",x"03",x"1b",
	x"28",x"a1",x"0f",x"05",x"24",x"31",x"0f",x"38",x"c9",x"ef",x"22",x"a3",x"03",x"1b",x"38",x"c9",
	x"ef",x"31",x"30",x"00",x"1e",x"a2",x"38",x"ef",x"01",x"31",x"30",x"00",x"07",x"25",x"04",x"38",
	x"c3",x"c4",x"36",x"02",x"31",x"30",x"00",x"09",x"a0",x"01",x"37",x"00",x"06",x"a1",x"01",x"05",
	x"02",x"a1",x"38",x"c9",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",
	x"10",x"10",x"10",x"00",x"10",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",
	x"7e",x"24",x"24",x"7e",x"24",x"00",x"00",x"08",x"3e",x"28",x"3e",x"0a",x"3e",x"08",x"00",x"62",
	x"64",x"08",x"10",x"26",x"46",x"00",x"00",x"10",x"28",x"10",x"2a",x"44",x"3a",x"00",x"00",x"08",
	x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"08",x"08",x"08",x"04",x"00",x"00",x"20",
	x"10",x"10",x"10",x"10",x"20",x"00",x"00",x"00",x"14",x"08",x"3e",x"08",x"14",x"00",x"00",x"00",
	x"08",x"08",x"3e",x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"10",x"00",x"00",
	x"00",x"00",x"3e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",
	x"02",x"04",x"08",x"10",x"20",x"00",x"00",x"3c",x"46",x"4a",x"52",x"62",x"3c",x"00",x"00",x"18",
	x"28",x"08",x"08",x"08",x"3e",x"00",x"00",x"3c",x"42",x"02",x"3c",x"40",x"7e",x"00",x"00",x"3c",
	x"42",x"0c",x"02",x"42",x"3c",x"00",x"00",x"08",x"18",x"28",x"48",x"7e",x"08",x"00",x"00",x"7e",
	x"40",x"7c",x"02",x"42",x"3c",x"00",x"00",x"3c",x"40",x"7c",x"42",x"42",x"3c",x"00",x"00",x"7e",
	x"02",x"04",x"08",x"10",x"10",x"00",x"00",x"3c",x"42",x"3c",x"42",x"42",x"3c",x"00",x"00",x"3c",
	x"42",x"42",x"3e",x"02",x"3c",x"00",x"00",x"00",x"00",x"10",x"00",x"00",x"10",x"00",x"00",x"00",
	x"10",x"00",x"00",x"10",x"10",x"20",x"00",x"00",x"04",x"08",x"10",x"08",x"04",x"00",x"00",x"00",
	x"00",x"3e",x"00",x"3e",x"00",x"00",x"00",x"00",x"10",x"08",x"04",x"08",x"10",x"00",x"00",x"3c",
	x"42",x"04",x"08",x"00",x"08",x"00",x"00",x"3c",x"4a",x"56",x"5e",x"40",x"3c",x"00",x"00",x"3c",
	x"42",x"42",x"7e",x"42",x"42",x"00",x"00",x"7c",x"42",x"7c",x"42",x"42",x"7c",x"00",x"00",x"3c",
	x"42",x"40",x"40",x"42",x"3c",x"00",x"00",x"78",x"44",x"42",x"42",x"44",x"78",x"00",x"00",x"7e",
	x"40",x"7c",x"40",x"40",x"7e",x"00",x"00",x"7e",x"40",x"7c",x"40",x"40",x"40",x"00",x"00",x"3c",
	x"42",x"40",x"4e",x"42",x"3c",x"00",x"00",x"42",x"42",x"7e",x"42",x"42",x"42",x"00",x"00",x"3e",
	x"08",x"08",x"08",x"08",x"3e",x"00",x"00",x"02",x"02",x"02",x"42",x"42",x"3c",x"00",x"00",x"44",
	x"48",x"70",x"48",x"44",x"42",x"00",x"00",x"40",x"40",x"40",x"40",x"40",x"7e",x"00",x"00",x"42",
	x"66",x"5a",x"42",x"42",x"42",x"00",x"00",x"42",x"62",x"52",x"4a",x"46",x"42",x"00",x"00",x"3c",
	x"42",x"42",x"42",x"42",x"3c",x"00",x"00",x"7c",x"42",x"42",x"7c",x"40",x"40",x"00",x"00",x"3c",
	x"42",x"42",x"52",x"4a",x"3c",x"00",x"00",x"7c",x"42",x"42",x"7c",x"44",x"42",x"00",x"00",x"3c",
	x"40",x"3c",x"02",x"42",x"3c",x"00",x"00",x"fe",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"42",
	x"42",x"42",x"42",x"42",x"3c",x"00",x"00",x"42",x"42",x"42",x"42",x"24",x"18",x"00",x"00",x"42",
	x"42",x"42",x"42",x"5a",x"24",x"00",x"00",x"42",x"24",x"18",x"18",x"24",x"42",x"00",x"00",x"82",
	x"44",x"28",x"10",x"10",x"10",x"00",x"00",x"7e",x"04",x"08",x"10",x"20",x"7e",x"00",x"00",x"0e",
	x"08",x"08",x"08",x"08",x"0e",x"00",x"00",x"00",x"40",x"20",x"10",x"08",x"04",x"00",x"00",x"70",
	x"10",x"10",x"10",x"10",x"70",x"00",x"00",x"10",x"38",x"54",x"10",x"10",x"10",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"ff",x"00",x"1c",x"22",x"78",x"20",x"20",x"7e",x"00",x"00",x"00",
	x"38",x"04",x"3c",x"44",x"3c",x"00",x"00",x"20",x"20",x"3c",x"22",x"22",x"3c",x"00",x"00",x"00",
	x"1c",x"20",x"20",x"20",x"1c",x"00",x"00",x"04",x"04",x"3c",x"44",x"44",x"3c",x"00",x"00",x"00",
	x"38",x"44",x"78",x"40",x"3c",x"00",x"00",x"0c",x"10",x"18",x"10",x"10",x"10",x"00",x"00",x"00",
	x"3c",x"44",x"44",x"3c",x"04",x"38",x"00",x"40",x"40",x"78",x"44",x"44",x"44",x"00",x"00",x"10",
	x"00",x"30",x"10",x"10",x"38",x"00",x"00",x"04",x"00",x"04",x"04",x"04",x"24",x"18",x"00",x"20",
	x"28",x"30",x"30",x"28",x"24",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"0c",x"00",x"00",x"00",
	x"68",x"54",x"54",x"54",x"54",x"00",x"00",x"00",x"78",x"44",x"44",x"44",x"44",x"00",x"00",x"00",
	x"38",x"44",x"44",x"44",x"38",x"00",x"00",x"00",x"78",x"44",x"44",x"78",x"40",x"40",x"00",x"00",
	x"3c",x"44",x"44",x"3c",x"04",x"06",x"00",x"00",x"1c",x"20",x"20",x"20",x"20",x"00",x"00",x"00",
	x"38",x"40",x"38",x"04",x"78",x"00",x"00",x"10",x"38",x"10",x"10",x"10",x"0c",x"00",x"00",x"00",
	x"44",x"44",x"44",x"44",x"38",x"00",x"00",x"00",x"44",x"44",x"28",x"28",x"10",x"00",x"00",x"00",
	x"44",x"54",x"54",x"54",x"28",x"00",x"00",x"00",x"44",x"28",x"10",x"28",x"44",x"00",x"00",x"00",
	x"44",x"44",x"44",x"3c",x"04",x"38",x"00",x"00",x"7c",x"08",x"10",x"20",x"7c",x"00",x"00",x"0e",
	x"08",x"30",x"08",x"08",x"0e",x"00",x"00",x"08",x"08",x"08",x"08",x"08",x"08",x"00",x"00",x"70",
	x"10",x"0c",x"10",x"10",x"70",x"00",x"00",x"14",x"28",x"00",x"00",x"00",x"00",x"00",x"3c",x"42",
	x"99",x"a1",x"a1",x"99",x"42",x"3c",

	others => x"07"
);

signal ReadAddress: std_logic_vector(Address'range);
signal DualReadAddress: std_logic_vector(DualAddress'range);

attribute syn_ramstyle: string;
attribute syn_ramstyle of RAM: signal is "block_ram";

begin

	process (Clock)
	begin
		if rising_edge(Clock) then
			if Enable = '1' and WriteEnable = '1' then
				RAM(conv_integer(Address)) <= DataIn;
			end if;

			if Enable = '1' then
				ReadAddress <= Address;
			end if;
			if DualEnable = '1' then
				DualReadAddress <= DualAddress;
			end if;
		end if;
	end process;

	DataOut <= RAM(conv_integer(ReadAddress));
	DualDataOut <= RAM(conv_integer(DualReadAddress));

end behavioral;
