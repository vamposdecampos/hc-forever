-- 32 Kbyte Block RAM, one R/W port, one read-only port

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity VideoRam is
generic (
	ADDR_BITS		: integer := 15;
	DATA_BITS		: integer := 8
);
port (
	Clock			: in  std_logic;
	Enable			: in  std_logic;
	WriteEnable		: in  std_logic;
	Address			: in  std_logic_vector(ADDR_BITS-1 downto 0);
	DataIn			: in  std_logic_vector(DATA_BITS-1 downto 0);
	DataOut			: out std_logic_vector(DATA_BITS-1 downto 0);

	DualEnable		: in  std_logic;
	DualAddress		: in  std_logic_vector(ADDR_BITS-1 downto 0);
	DualDataOut		: out std_logic_vector(DATA_BITS-1 downto 0)
);
end VideoRam;

architecture behavioral of VideoRam is

type ram_type is array (0 to 2**ADDR_BITS - 1) of std_logic_vector (DataOut'range);
signal RAM: ram_type := (

	x"f3",x"3e",x"3f",x"ed",x"47",x"31",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"21",x"3a",
	x"01",x"22",x"1a",x"60",x"cd",x"1a",x"00",x"c3",x"75",x"05",x"cd",x"18",x"02",x"06",x"1a",x"21",
	x"00",x"60",x"36",x"00",x"23",x"10",x"fb",x"21",x"d7",x"0a",x"22",x"00",x"60",x"3e",x"06",x"32",
	x"02",x"60",x"cd",x"f0",x"00",x"21",x"b4",x"2d",x"22",x"00",x"60",x"3e",x"1e",x"32",x"02",x"60",
	x"cd",x"f0",x"00",x"3e",x"19",x"32",x"02",x"60",x"cd",x"41",x"01",x"3e",x"1f",x"32",x"02",x"60",
	x"cd",x"41",x"01",x"3e",x"26",x"32",x"02",x"60",x"cd",x"41",x"01",x"3e",x"0c",x"32",x"9b",x"6e",
	x"af",x"32",x"9c",x"6e",x"3e",x"08",x"32",x"a1",x"6e",x"3e",x"02",x"32",x"9f",x"6e",x"32",x"a0",
	x"6e",x"21",x"c9",x"00",x"22",x"a2",x"6e",x"2a",x"e6",x"00",x"22",x"9d",x"6e",x"cd",x"a1",x"17",
	x"21",x"cf",x"00",x"22",x"a2",x"6e",x"2a",x"e8",x"00",x"22",x"9d",x"6e",x"cd",x"a1",x"17",x"3e",
	x"08",x"32",x"a1",x"6e",x"3e",x"04",x"32",x"9f",x"6e",x"32",x"a0",x"6e",x"21",x"d8",x"00",x"22",
	x"a2",x"6e",x"2a",x"ea",x"00",x"22",x"9d",x"6e",x"cd",x"a1",x"17",x"21",x"de",x"00",x"22",x"a2",
	x"6e",x"2a",x"ec",x"00",x"22",x"9d",x"6e",x"cd",x"a1",x"17",x"06",x"0a",x"c5",x"01",x"ff",x"ff",
	x"0d",x"20",x"fd",x"10",x"fb",x"c1",x"10",x"f4",x"c9",x"50",x"53",x"49",x"4f",x"4e",x"ff",x"53",
	x"4f",x"46",x"54",x"57",x"41",x"52",x"45",x"ff",x"53",x"50",x"41",x"43",x"45",x"ff",x"52",x"41",
	x"49",x"44",x"45",x"52",x"53",x"ff",x"19",x"23",x"05",x"32",x"2a",x"64",x"16",x"87",x"c8",x"03",
	x"af",x"cd",x"6a",x"13",x"21",x"00",x"03",x"22",x"04",x"60",x"2a",x"04",x"60",x"cd",x"67",x"17",
	x"ed",x"5b",x"02",x"60",x"cd",x"82",x"13",x"22",x"06",x"60",x"2a",x"04",x"60",x"cd",x"9c",x"17",
	x"ed",x"5b",x"02",x"60",x"cd",x"82",x"13",x"3a",x"00",x"60",x"85",x"4f",x"3a",x"00",x"60",x"95",
	x"6f",x"3a",x"06",x"60",x"47",x"3a",x"01",x"60",x"80",x"47",x"60",x"cd",x"ec",x"12",x"ed",x"4b",
	x"04",x"60",x"0b",x"0b",x"ed",x"43",x"04",x"60",x"21",x"00",x"01",x"b7",x"ed",x"42",x"38",x"ba",
	x"c9",x"21",x"00",x"04",x"22",x"04",x"60",x"3a",x"02",x"60",x"cb",x"3f",x"32",x"0a",x"60",x"3a",
	x"02",x"60",x"cb",x"27",x"32",x"08",x"60",x"2a",x"ee",x"00",x"cd",x"67",x"17",x"32",x"0c",x"60",
	x"ed",x"5b",x"08",x"60",x"cd",x"82",x"13",x"22",x"0e",x"60",x"3a",x"0c",x"60",x"ed",x"5b",x"0a",
	x"60",x"cd",x"82",x"13",x"22",x"10",x"60",x"2a",x"ee",x"00",x"cd",x"9c",x"17",x"32",x"0d",x"60",
	x"ed",x"5b",x"08",x"60",x"cd",x"82",x"13",x"22",x"12",x"60",x"ed",x"5b",x"0a",x"60",x"3a",x"0d",
	x"60",x"cd",x"82",x"13",x"22",x"14",x"60",x"2a",x"04",x"60",x"cd",x"9c",x"17",x"ed",x"5b",x"12",
	x"60",x"cd",x"82",x"13",x"22",x"16",x"60",x"2a",x"04",x"60",x"cd",x"67",x"17",x"ed",x"5b",x"10",
	x"60",x"cd",x"82",x"13",x"ed",x"4b",x"16",x"60",x"09",x"3a",x"00",x"60",x"85",x"32",x"16",x"60",
	x"2a",x"04",x"60",x"cd",x"67",x"17",x"ed",x"5b",x"14",x"60",x"cd",x"82",x"13",x"22",x"18",x"60",
	x"2a",x"04",x"60",x"cd",x"9c",x"17",x"ed",x"5b",x"0e",x"60",x"cd",x"82",x"13",x"ed",x"5b",x"18",
	x"60",x"eb",x"b7",x"ed",x"52",x"3a",x"01",x"60",x"85",x"47",x"3a",x"16",x"60",x"4f",x"ed",x"5b",
	x"04",x"60",x"b7",x"21",x"fe",x"01",x"ed",x"52",x"30",x"05",x"cd",x"42",x"14",x"18",x"03",x"cd",
	x"4f",x"14",x"ed",x"4b",x"04",x"60",x"0b",x"0b",x"0b",x"0b",x"ed",x"43",x"04",x"60",x"21",x"00",
	x"00",x"b7",x"ed",x"42",x"da",x"97",x"01",x"c9",x"cd",x"ad",x"12",x"3e",x"01",x"32",x"48",x"5c",
	x"3e",x"01",x"d3",x"fe",x"3e",x"0e",x"57",x"5f",x"21",x"00",x"00",x"39",x"31",x"00",x"5b",x"01",
	x"80",x"01",x"d5",x"0b",x"79",x"b0",x"20",x"fa",x"f9",x"c9",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"00",x"10",x"00",x"00",x"24",x"24",x"00",x"00",x"00",
	x"00",x"00",x"00",x"24",x"7e",x"24",x"24",x"7e",x"24",x"00",x"00",x"08",x"3e",x"28",x"3e",x"0a",
	x"3e",x"08",x"00",x"62",x"64",x"08",x"10",x"26",x"46",x"00",x"00",x"10",x"28",x"10",x"2a",x"44",
	x"3a",x"00",x"00",x"08",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"08",x"08",x"08",
	x"04",x"00",x"00",x"20",x"10",x"10",x"10",x"10",x"20",x"00",x"00",x"00",x"14",x"08",x"3e",x"08",
	x"14",x"00",x"00",x"00",x"08",x"08",x"3e",x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"08",
	x"08",x"10",x"00",x"00",x"00",x"00",x"3e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",
	x"18",x"00",x"00",x"00",x"02",x"04",x"08",x"10",x"20",x"00",x"00",x"3c",x"46",x"4a",x"52",x"62",
	x"3c",x"00",x"00",x"18",x"28",x"08",x"08",x"08",x"3e",x"00",x"00",x"3c",x"42",x"02",x"3c",x"40",
	x"7e",x"00",x"00",x"3c",x"42",x"0c",x"02",x"42",x"3c",x"00",x"00",x"08",x"18",x"28",x"48",x"7e",
	x"08",x"00",x"00",x"7e",x"40",x"7c",x"02",x"42",x"3c",x"00",x"00",x"3c",x"40",x"7c",x"42",x"42",
	x"3c",x"00",x"00",x"7e",x"02",x"04",x"08",x"10",x"10",x"00",x"00",x"3c",x"42",x"3c",x"42",x"42",
	x"3c",x"00",x"00",x"3c",x"42",x"42",x"3e",x"02",x"3c",x"00",x"00",x"00",x"00",x"10",x"00",x"00",
	x"10",x"00",x"00",x"00",x"10",x"00",x"00",x"10",x"10",x"20",x"00",x"00",x"04",x"08",x"10",x"08",
	x"04",x"00",x"00",x"00",x"00",x"3e",x"00",x"3e",x"00",x"00",x"00",x"00",x"10",x"08",x"04",x"08",
	x"10",x"00",x"00",x"3c",x"42",x"04",x"08",x"00",x"08",x"00",x"00",x"3c",x"4a",x"56",x"5e",x"40",
	x"3c",x"00",x"00",x"3c",x"42",x"42",x"7e",x"42",x"42",x"00",x"00",x"7c",x"42",x"7c",x"42",x"42",
	x"7c",x"00",x"00",x"3c",x"42",x"40",x"40",x"42",x"3c",x"00",x"00",x"78",x"44",x"42",x"42",x"44",
	x"78",x"00",x"00",x"7e",x"40",x"7c",x"40",x"40",x"7e",x"00",x"00",x"7e",x"40",x"7c",x"40",x"40",
	x"40",x"00",x"00",x"3c",x"42",x"40",x"4e",x"42",x"3c",x"00",x"00",x"42",x"42",x"7e",x"42",x"42",
	x"42",x"00",x"00",x"3e",x"08",x"08",x"08",x"08",x"3e",x"00",x"00",x"02",x"02",x"02",x"42",x"42",
	x"3c",x"00",x"00",x"44",x"48",x"70",x"48",x"44",x"42",x"00",x"00",x"40",x"40",x"40",x"40",x"40",
	x"7e",x"00",x"00",x"42",x"66",x"5a",x"42",x"42",x"42",x"00",x"00",x"42",x"62",x"52",x"4a",x"46",
	x"42",x"00",x"00",x"3c",x"42",x"42",x"42",x"42",x"3c",x"00",x"00",x"7c",x"42",x"42",x"7c",x"40",
	x"40",x"00",x"00",x"3c",x"42",x"42",x"52",x"4a",x"3c",x"00",x"00",x"7c",x"42",x"42",x"7c",x"44",
	x"42",x"00",x"00",x"3c",x"40",x"3c",x"02",x"42",x"3c",x"00",x"00",x"fe",x"10",x"10",x"10",x"10",
	x"10",x"00",x"00",x"42",x"42",x"42",x"42",x"42",x"3c",x"00",x"00",x"42",x"42",x"42",x"42",x"24",
	x"18",x"00",x"00",x"42",x"42",x"42",x"42",x"5a",x"24",x"00",x"00",x"42",x"24",x"18",x"18",x"24",
	x"42",x"00",x"00",x"82",x"44",x"28",x"10",x"10",x"10",x"00",x"00",x"7e",x"04",x"08",x"10",x"20",
	x"7e",x"00",x"00",x"0e",x"08",x"08",x"08",x"08",x"0e",x"00",x"00",x"00",x"40",x"20",x"10",x"08",
	x"04",x"00",x"00",x"70",x"10",x"10",x"10",x"10",x"70",x"00",x"00",x"10",x"38",x"54",x"10",x"10",
	x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"ff",x"00",x"1c",x"22",x"78",x"20",x"20",
	x"7e",x"00",x"00",x"00",x"38",x"04",x"3c",x"44",x"3c",x"00",x"00",x"20",x"20",x"3c",x"22",x"22",
	x"3c",x"00",x"00",x"00",x"1c",x"20",x"20",x"20",x"1c",x"00",x"00",x"04",x"04",x"3c",x"44",x"44",
	x"3c",x"00",x"00",x"00",x"38",x"44",x"78",x"40",x"3c",x"00",x"00",x"0c",x"10",x"18",x"10",x"10",
	x"10",x"00",x"00",x"00",x"3c",x"44",x"44",x"3c",x"04",x"38",x"00",x"40",x"40",x"78",x"44",x"44",
	x"44",x"00",x"00",x"10",x"00",x"30",x"10",x"10",x"38",x"00",x"00",x"04",x"00",x"04",x"04",x"04",
	x"24",x"18",x"00",x"20",x"28",x"30",x"30",x"28",x"24",x"00",x"00",x"10",x"10",x"10",x"10",x"10",
	x"0c",x"00",x"00",x"00",x"68",x"54",x"54",x"54",x"54",x"00",x"00",x"00",x"78",x"44",x"44",x"44",
	x"44",x"00",x"00",x"00",x"38",x"44",x"44",x"44",x"38",x"00",x"00",x"00",x"78",x"44",x"44",x"78",
	x"40",x"40",x"00",x"00",x"3c",x"44",x"44",x"3c",x"04",x"06",x"00",x"00",x"1c",x"20",x"20",x"20",
	x"20",x"00",x"00",x"00",x"38",x"40",x"38",x"04",x"78",x"00",x"00",x"10",x"38",x"10",x"10",x"10",
	x"0c",x"00",x"00",x"00",x"44",x"44",x"44",x"44",x"38",x"00",x"00",x"00",x"44",x"44",x"28",x"28",
	x"10",x"00",x"00",x"00",x"44",x"54",x"54",x"54",x"28",x"00",x"00",x"00",x"44",x"28",x"10",x"28",
	x"44",x"00",x"00",x"00",x"44",x"44",x"44",x"3c",x"04",x"38",x"00",x"00",x"7c",x"08",x"10",x"20",
	x"7c",x"00",x"00",x"0e",x"08",x"30",x"08",x"08",x"0e",x"00",x"00",x"08",x"08",x"08",x"08",x"08",
	x"08",x"00",x"00",x"70",x"10",x"0c",x"10",x"10",x"70",x"00",x"00",x"14",x"28",x"00",x"00",x"00",
	x"00",x"00",x"3c",x"42",x"99",x"a1",x"a1",x"99",x"42",x"3c",x"05",x"06",x"04",x"04",x"02",x"02",
	x"07",x"03",x"01",x"01",x"01",x"00",x"00",x"00",x"03",x"05",x"00",x"00",x"37",x"0b",x"0b",x"0b",
	x"0b",x"0b",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"00",x"00",x"04",
	x"01",x"00",x"0b",x"00",x"b8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"08",x"f3",x"31",x"00",x"80",x"21",x"00",x"00",x"22",x"1e",x"60",x"22",
	x"1c",x"60",x"21",x"35",x"82",x"22",x"a4",x"6e",x"22",x"a6",x"6e",x"cd",x"01",x"06",x"cd",x"ad",
	x"12",x"cd",x"ab",x"06",x"cd",x"d7",x"06",x"cd",x"12",x"06",x"cd",x"f0",x"05",x"cd",x"8e",x"0e",
	x"cd",x"99",x"07",x"cd",x"4e",x"0e",x"cd",x"e9",x"11",x"cd",x"8e",x"10",x"cd",x"1e",x"07",x"cd",
	x"13",x"07",x"cd",x"c1",x"0c",x"cd",x"bb",x"0a",x"3a",x"2a",x"60",x"b7",x"ca",x"66",x"06",x"cd",
	x"71",x"09",x"28",x"0a",x"3a",x"26",x"60",x"b7",x"ca",x"55",x"07",x"cd",x"d7",x"06",x"cd",x"6b",
	x"08",x"cd",x"e5",x"05",x"3a",x"26",x"60",x"b7",x"ca",x"55",x"07",x"3a",x"28",x"60",x"b7",x"c2",
	x"55",x"07",x"c3",x"33",x"06",x"3a",x"53",x"60",x"3d",x"32",x"53",x"60",x"c0",x"cd",x"b4",x"0f",
	x"3a",x"2a",x"60",x"cb",x"3f",x"cb",x"3f",x"47",x"cb",x"3f",x"80",x"c6",x"04",x"32",x"53",x"60",
	x"c9",x"3e",x"01",x"32",x"56",x"60",x"21",x"42",x"05",x"11",x"20",x"60",x"01",x"0a",x"00",x"ed",
	x"b0",x"c9",x"21",x"4c",x"05",x"11",x"2a",x"60",x"01",x"29",x"00",x"ed",x"b0",x"3a",x"23",x"60",
	x"3c",x"c8",x"32",x"23",x"60",x"fe",x"32",x"d0",x"fe",x"09",x"d8",x"3a",x"27",x"60",x"3c",x"32",
	x"27",x"60",x"c9",x"3a",x"50",x"60",x"b7",x"20",x"06",x"3a",x"20",x"60",x"cd",x"5b",x"06",x"3a",
	x"43",x"60",x"b7",x"20",x"06",x"3a",x"21",x"60",x"cd",x"5b",x"06",x"3a",x"44",x"60",x"b7",x"c2",
	x"ac",x"05",x"3a",x"22",x"60",x"cd",x"5b",x"06",x"c3",x"ac",x"05",x"47",x"c5",x"06",x"00",x"00",
	x"10",x"fd",x"c1",x"10",x"f7",x"c9",x"3a",x"29",x"60",x"3c",x"fe",x"08",x"20",x"01",x"3d",x"32",
	x"29",x"60",x"c3",x"97",x"05",x"32",x"54",x"60",x"c5",x"cd",x"c6",x"12",x"3a",x"54",x"60",x"ed",
	x"44",x"c6",x"05",x"28",x"05",x"dd",x"23",x"3d",x"20",x"fb",x"dd",x"7e",x"00",x"dd",x"23",x"cd",
	x"cb",x"13",x"c1",x"50",x"59",x"1c",x"d5",x"cd",x"52",x"13",x"3a",x"54",x"60",x"3d",x"32",x"54",
	x"60",x"20",x"e7",x"af",x"cd",x"cb",x"13",x"c1",x"c3",x"52",x"13",x"ed",x"5b",x"1c",x"60",x"2a",
	x"1e",x"60",x"b7",x"ed",x"52",x"30",x"04",x"ed",x"53",x"1e",x"60",x"21",x"00",x"00",x"22",x"1c",
	x"60",x"cd",x"88",x"15",x"15",x"00",x"48",x"49",x"47",x"48",x"20",x"00",x"01",x"1a",x"00",x"2a",
	x"1e",x"60",x"3e",x"05",x"c3",x"75",x"06",x"11",x"00",x"40",x"cd",x"99",x"0a",x"3a",x"26",x"60",
	x"3d",x"28",x"2d",x"fa",x"10",x"07",x"32",x"55",x"60",x"ed",x"5b",x"41",x"60",x"d5",x"af",x"32",
	x"42",x"60",x"3e",x"48",x"32",x"41",x"60",x"cd",x"4e",x"0e",x"3a",x"41",x"60",x"c6",x"18",x"32",
	x"41",x"60",x"3a",x"55",x"60",x"3d",x"32",x"55",x"60",x"20",x"ec",x"d1",x"ed",x"53",x"41",x"60",
	x"cd",x"c1",x"06",x"2a",x"1c",x"60",x"01",x"00",x"00",x"3e",x"05",x"c3",x"75",x"06",x"3a",x"24",
	x"60",x"b7",x"c0",x"2a",x"1c",x"60",x"01",x"64",x"00",x"ed",x"42",x"d8",x"3e",x"01",x"32",x"24",
	x"60",x"3a",x"26",x"60",x"3c",x"32",x"26",x"60",x"06",x"08",x"3a",x"48",x"5c",x"c6",x"08",x"e6",
	x"38",x"32",x"48",x"5c",x"cd",x"0d",x"16",x"0c",x"28",x"12",x"1e",x"18",x"14",x"30",x"0a",x"00",
	x"10",x"e8",x"c3",x"d7",x"06",x"cd",x"88",x"15",x"00",x"17",x"47",x"41",x"4d",x"45",x"20",x"4f",
	x"56",x"45",x"52",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"48",x"49",x"54",x"20",x"46",x"49",
	x"52",x"45",x"20",x"54",x"4f",x"20",x"50",x"4c",x"41",x"59",x"00",x"06",x"19",x"cd",x"0d",x"16",
	x"28",x"32",x"28",x"28",x"28",x"1e",x"28",x"14",x"28",x"0a",x"00",x"10",x"f0",x"cd",x"d6",x"0c",
	x"3a",x"4f",x"60",x"b7",x"28",x"f7",x"c3",x"8b",x"05",x"3a",x"3a",x"05",x"e6",x"38",x"32",x"48",
	x"5c",x"3a",x"3a",x"05",x"01",x"03",x"00",x"21",x"00",x"58",x"77",x"23",x"10",x"fc",x"0d",x"20",
	x"f9",x"cd",x"0d",x"16",x"64",x"64",x"00",x"01",x"00",x"01",x"3a",x"41",x"05",x"5f",x"16",x"20",
	x"cd",x"59",x"11",x"01",x"00",x"17",x"3a",x"40",x"05",x"5f",x"16",x"20",x"c3",x"59",x"11",x"13",
	x"01",x"14",x"02",x"03",x"03",x"07",x"03",x"0c",x"03",x"11",x"03",x"15",x"03",x"02",x"04",x"07",
	x"04",x"0c",x"04",x"11",x"04",x"16",x"04",x"03",x"05",x"07",x"05",x"0c",x"05",x"11",x"05",x"15",
	x"05",x"14",x"06",x"13",x"07",x"ff",x"03",x"01",x"02",x"02",x"01",x"03",x"05",x"03",x"0a",x"03",
	x"0f",x"03",x"13",x"03",x"00",x"04",x"05",x"04",x"0a",x"04",x"0f",x"04",x"14",x"04",x"01",x"05",
	x"05",x"05",x"0a",x"05",x"0f",x"05",x"13",x"05",x"02",x"06",x"03",x"07",x"ff",x"04",x"01",x"03",
	x"02",x"02",x"03",x"06",x"03",x"0b",x"03",x"10",x"03",x"14",x"03",x"01",x"04",x"06",x"04",x"0b",
	x"04",x"10",x"04",x"15",x"04",x"02",x"05",x"06",x"05",x"0b",x"05",x"10",x"05",x"14",x"05",x"03",
	x"06",x"04",x"07",x"ff",x"14",x"01",x"15",x"02",x"04",x"03",x"08",x"03",x"0d",x"03",x"12",x"03",
	x"16",x"03",x"03",x"04",x"08",x"04",x"0d",x"04",x"12",x"04",x"17",x"04",x"04",x"05",x"08",x"05",
	x"0d",x"05",x"12",x"05",x"16",x"05",x"15",x"06",x"14",x"07",x"ff",x"3a",x"50",x"60",x"b7",x"20",
	x"28",x"3a",x"a6",x"6e",x"fe",x"ff",x"c0",x"3a",x"a7",x"6e",x"fe",x"19",x"d0",x"3a",x"a7",x"6e",
	x"cb",x"47",x"28",x"0a",x"3e",x"01",x"32",x"50",x"60",x"af",x"32",x"51",x"60",x"c9",x"3e",x"ff",
	x"32",x"50",x"60",x"3e",x"e9",x"32",x"51",x"60",x"c9",x"3a",x"56",x"60",x"ed",x"44",x"32",x"56",
	x"60",x"f2",x"25",x"09",x"dd",x"21",x"51",x"60",x"3a",x"50",x"60",x"fe",x"01",x"28",x"0e",x"21",
	x"cf",x"07",x"dd",x"35",x"00",x"af",x"dd",x"be",x"00",x"20",x"19",x"18",x"0d",x"21",x"1d",x"08",
	x"dd",x"34",x"00",x"3e",x"ea",x"dd",x"be",x"00",x"20",x"0a",x"af",x"32",x"50",x"60",x"11",x"20",
	x"40",x"c3",x"99",x"0a",x"3e",x"01",x"cd",x"2a",x"14",x"af",x"cd",x"2a",x"14",x"3a",x"44",x"60",
	x"b7",x"c8",x"dd",x"21",x"45",x"60",x"dd",x"7e",x"01",x"fe",x"10",x"d0",x"3a",x"51",x"60",x"dd",
	x"be",x"00",x"d0",x"c6",x"17",x"dd",x"be",x"00",x"d8",x"cd",x"01",x"09",x"af",x"32",x"50",x"60",
	x"c9",x"cd",x"ca",x"08",x"cd",x"34",x"09",x"cd",x"0d",x"16",x"0a",x"ff",x"0a",x"c8",x"14",x"96",
	x"05",x"c8",x"14",x"96",x"14",x"78",x"14",x"64",x"14",x"50",x"14",x"3c",x"14",x"28",x"00",x"11",
	x"20",x"40",x"c3",x"99",x"0a",x"cd",x"0d",x"16",x"02",x"19",x"02",x"32",x"02",x"19",x"00",x"c9",
	x"05",x"05",x"0a",x"14",x"3a",x"a7",x"6e",x"1f",x"e6",x"03",x"21",x"30",x"09",x"cd",x"5f",x"09",
	x"7e",x"47",x"2a",x"1c",x"60",x"cd",x"5f",x"09",x"22",x"1c",x"60",x"3a",x"51",x"60",x"cb",x"3f",
	x"cb",x"3f",x"cb",x"3f",x"4f",x"68",x"26",x"00",x"06",x"01",x"3e",x"02",x"c3",x"75",x"06",x"85",
	x"6f",x"d0",x"24",x"c9",x"00",x"00",x"00",x"01",x"00",x"02",x"00",x"03",x"00",x"04",x"00",x"05",
	x"ff",x"3e",x"04",x"32",x"5a",x"60",x"dd",x"21",x"47",x"60",x"dd",x"7e",x"01",x"b7",x"28",x"05",
	x"cd",x"02",x"0a",x"18",x"03",x"cd",x"9a",x"09",x"cd",x"8e",x"09",x"20",x"ed",x"c9",x"dd",x"23",
	x"dd",x"23",x"3a",x"5a",x"60",x"3d",x"32",x"5a",x"60",x"c9",x"cd",x"b6",x"18",x"3a",x"a4",x"6e",
	x"47",x"3a",x"27",x"60",x"b7",x"c8",x"b8",x"d8",x"3a",x"3d",x"60",x"32",x"57",x"60",x"3a",x"41",
	x"60",x"c6",x"07",x"47",x"3a",x"a6",x"6e",x"e6",x"0f",x"80",x"32",x"58",x"60",x"3a",x"a5",x"6e",
	x"fe",x"7f",x"30",x"06",x"3a",x"a6",x"6e",x"32",x"58",x"60",x"3a",x"57",x"60",x"dd",x"e5",x"cd",
	x"d1",x"0e",x"dd",x"7e",x"01",x"32",x"59",x"60",x"3a",x"58",x"60",x"cd",x"26",x"0b",x"dd",x"e1",
	x"20",x"0b",x"3a",x"57",x"60",x"3d",x"32",x"57",x"60",x"f2",x"ca",x"09",x"c9",x"3a",x"59",x"60",
	x"3c",x"3c",x"cb",x"27",x"cb",x"27",x"cb",x"27",x"dd",x"77",x"01",x"3a",x"58",x"60",x"dd",x"77",
	x"00",x"c9",x"21",x"64",x"09",x"3e",x"01",x"cd",x"2a",x"14",x"dd",x"7e",x"01",x"3c",x"fe",x"b9",
	x"d2",x"b6",x"0a",x"fe",x"b1",x"d2",x"32",x"0a",x"dd",x"77",x"01",x"c6",x"05",x"47",x"dd",x"4e",
	x"00",x"dd",x"e5",x"cd",x"42",x"12",x"dd",x"e1",x"c2",x"b6",x"0a",x"21",x"64",x"09",x"af",x"c3",
	x"2a",x"14",x"dd",x"7e",x"00",x"47",x"3a",x"41",x"60",x"b8",x"30",x"53",x"c6",x"13",x"b8",x"38",
	x"4e",x"af",x"32",x"41",x"60",x"06",x"08",x"3a",x"48",x"5c",x"c6",x"08",x"e6",x"38",x"32",x"48",
	x"5c",x"cd",x"0d",x"16",x"28",x"0a",x"28",x"14",x"28",x"28",x"28",x"50",x"00",x"10",x"e8",x"cd",
	x"96",x"0a",x"cd",x"0d",x"16",x"32",x"ff",x"ff",x"32",x"32",x"ff",x"00",x"3a",x"26",x"60",x"3d",
	x"32",x"26",x"60",x"c4",x"4e",x"0e",x"cd",x"7d",x"0a",x"f6",x"01",x"e1",x"c9",x"3e",x"04",x"32",
	x"5a",x"60",x"dd",x"21",x"47",x"60",x"cd",x"a9",x"0a",x"cd",x"8e",x"09",x"20",x"f8",x"c9",x"dd",
	x"7e",x"01",x"3c",x"c3",x"18",x"0a",x"11",x"e0",x"50",x"0e",x"08",x"af",x"06",x"20",x"d5",x"12",
	x"13",x"10",x"fc",x"d1",x"14",x"0d",x"20",x"f4",x"c9",x"dd",x"7e",x"01",x"b7",x"c8",x"21",x"64",
	x"09",x"3e",x"01",x"cd",x"2a",x"14",x"dd",x"36",x"01",x"00",x"c9",x"3a",x"44",x"60",x"b7",x"c8",
	x"cd",x"c6",x"0a",x"c3",x"75",x"0c",x"3a",x"46",x"60",x"cb",x"3f",x"cb",x"3f",x"cb",x"3f",x"3c",
	x"32",x"5f",x"60",x"3a",x"3d",x"60",x"32",x"5d",x"60",x"cd",x"d1",x"0e",x"3a",x"5f",x"60",x"dd",
	x"be",x"01",x"28",x"08",x"3a",x"5d",x"60",x"3d",x"f2",x"d6",x"0a",x"c9",x"3a",x"45",x"60",x"cd",
	x"26",x"0b",x"c8",x"c3",x"6d",x"0b",x"10",x"80",x"09",x"10",x"49",x"20",x"26",x"40",x"10",x"80",
	x"00",x"00",x"10",x"80",x"66",x"60",x"89",x"30",x"09",x"80",x"10",x"80",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"32",x"5b",x"60",x"cd",x"ae",x"10",x"dd",x"21",x"35",x"6e",
	x"3a",x"5b",x"60",x"47",x"cb",x"3f",x"cb",x"3f",x"cb",x"3f",x"32",x"5e",x"60",x"dd",x"96",x"04",
	x"38",x"29",x"cb",x"47",x"28",x"04",x"cb",x"50",x"20",x"21",x"dd",x"be",x"05",x"30",x"1c",x"e6",
	x"fe",x"dd",x"86",x"04",x"32",x"5e",x"60",x"dd",x"96",x"02",x"32",x"5c",x"60",x"4f",x"06",x"00",
	x"dd",x"2a",x"35",x"6e",x"dd",x"09",x"dd",x"7e",x"02",x"b7",x"c9",x"af",x"c9",x"cd",x"cc",x"0b",
	x"21",x"f6",x"0a",x"22",x"60",x"60",x"21",x"06",x"0b",x"22",x"62",x"60",x"cd",x"dd",x"0b",x"cd",
	x"3d",x"0e",x"cd",x"0d",x"16",x"10",x"50",x"20",x"28",x"40",x"14",x"80",x"0a",x"00",x"cd",x"5c",
	x"0c",x"21",x"16",x"0b",x"22",x"60",x"60",x"22",x"62",x"60",x"cd",x"dd",x"0b",x"3a",x"2a",x"60",
	x"3d",x"32",x"2a",x"60",x"c2",x"03",x"0c",x"cd",x"7d",x"0a",x"06",x"28",x"3a",x"48",x"5c",x"c6",
	x"08",x"e6",x"38",x"32",x"48",x"5c",x"cd",x"0d",x"16",x"10",x"64",x"20",x"32",x"40",x"19",x"20",
	x"32",x"00",x"10",x"e8",x"cd",x"ca",x"08",x"cd",x"96",x"0a",x"e1",x"c9",x"06",x"20",x"11",x"16",
	x"00",x"af",x"dd",x"77",x"02",x"dd",x"77",x"03",x"dd",x"19",x"10",x"f6",x"c9",x"ed",x"4b",x"5e",
	x"60",x"cd",x"f8",x"15",x"2a",x"60",x"60",x"cd",x"f5",x"0b",x"ed",x"4b",x"5e",x"60",x"04",x"cd",
	x"f8",x"15",x"2a",x"62",x"60",x"06",x"08",x"ed",x"a0",x"ed",x"a0",x"1b",x"1b",x"03",x"03",x"14",
	x"10",x"f5",x"c9",x"21",x"2b",x"60",x"3a",x"5d",x"60",x"cd",x"70",x"0c",x"35",x"21",x"30",x"60",
	x"dd",x"21",x"35",x"6e",x"3a",x"5c",x"60",x"cb",x"3f",x"cd",x"70",x"0c",x"35",x"21",x"2b",x"60",
	x"3a",x"3d",x"60",x"3c",x"47",x"cd",x"70",x"0c",x"af",x"2b",x"05",x"b6",x"28",x"fb",x"78",x"32",
	x"3d",x"60",x"06",x"ff",x"21",x"30",x"60",x"af",x"2b",x"23",x"04",x"b6",x"28",x"fb",x"78",x"32",
	x"3f",x"60",x"21",x"30",x"60",x"3e",x"0b",x"47",x"04",x"cd",x"70",x"0c",x"af",x"2b",x"05",x"b6",
	x"28",x"fb",x"78",x"32",x"40",x"60",x"c9",x"03",x"02",x"02",x"01",x"01",x"3a",x"5d",x"60",x"21",
	x"57",x"0c",x"cd",x"70",x"0c",x"7e",x"2a",x"1c",x"60",x"cd",x"70",x"0c",x"22",x"1c",x"60",x"c9",
	x"85",x"6f",x"d0",x"24",x"c9",x"dd",x"21",x"47",x"60",x"3e",x"04",x"32",x"64",x"60",x"ed",x"4b",
	x"45",x"60",x"dd",x"7e",x"01",x"b7",x"28",x"20",x"dd",x"7e",x"00",x"b9",x"20",x"1a",x"dd",x"7e",
	x"01",x"90",x"ed",x"44",x"fe",x"06",x"30",x"10",x"cd",x"a9",x"0a",x"cd",x"0d",x"16",x"04",x"18",
	x"08",x"0c",x"10",x"06",x"00",x"c3",x"3d",x"0e",x"dd",x"23",x"dd",x"23",x"3a",x"64",x"60",x"3d",
	x"32",x"64",x"60",x"20",x"cd",x"ed",x"4b",x"45",x"60",x"05",x"cd",x"42",x"12",x"c8",x"c3",x"3d",
	x"0e",x"cd",x"d6",x"0c",x"cd",x"2e",x"0d",x"3a",x"44",x"60",x"b7",x"c2",x"1e",x"0e",x"3a",x"4f",
	x"60",x"b7",x"c8",x"c3",x"fd",x"0d",x"01",x"fe",x"fe",x"ed",x"58",x"01",x"fe",x"f7",x"ed",x"50",
	x"3a",x"41",x"60",x"0e",x"00",x"cb",x"4b",x"28",x"04",x"cb",x"42",x"20",x"04",x"b7",x"28",x"01",
	x"0d",x"cb",x"53",x"28",x"04",x"cb",x"4a",x"20",x"05",x"fe",x"eb",x"28",x"01",x"0c",x"79",x"32",
	x"43",x"60",x"01",x"fe",x"7f",x"ed",x"58",x"cb",x"43",x"28",x"0e",x"cb",x"62",x"28",x"0a",x"3e",
	x"01",x"32",x"65",x"60",x"af",x"32",x"4f",x"60",x"c9",x"cb",x"63",x"20",x"02",x"c1",x"c9",x"3a",
	x"65",x"60",x"b7",x"ca",x"14",x"0d",x"32",x"4f",x"60",x"af",x"32",x"65",x"60",x"c9",x"3a",x"43",
	x"60",x"b7",x"c8",x"f2",x"37",x"0d",x"af",x"dd",x"21",x"41",x"60",x"cd",x"53",x"0d",x"3e",x"01",
	x"cd",x"2a",x"14",x"af",x"cd",x"2a",x"14",x"3a",x"43",x"60",x"47",x"3a",x"41",x"60",x"80",x"32",
	x"41",x"60",x"c9",x"21",x"5c",x"0d",x"b7",x"c0",x"21",x"a6",x"0d",x"c9",x"0a",x"00",x"09",x"01",
	x"01",x"02",x"09",x"02",x"13",x"02",x"01",x"03",x"09",x"03",x"13",x"03",x"01",x"04",x"06",x"04",
	x"12",x"04",x"01",x"05",x"01",x"06",x"06",x"06",x"12",x"06",x"01",x"07",x"07",x"07",x"13",x"07",
	x"ff",x"0b",x"00",x"0c",x"01",x"02",x"02",x"0c",x"02",x"14",x"02",x"02",x"03",x"0c",x"03",x"14",
	x"03",x"03",x"04",x"0f",x"04",x"14",x"04",x"14",x"05",x"03",x"06",x"0f",x"06",x"14",x"06",x"02",
	x"07",x"0e",x"07",x"14",x"07",x"ff",x"0a",x"00",x"0b",x"01",x"01",x"02",x"0b",x"02",x"13",x"02",
	x"01",x"03",x"0b",x"03",x"13",x"03",x"02",x"04",x"0e",x"04",x"13",x"04",x"13",x"05",x"02",x"06",
	x"0e",x"06",x"13",x"06",x"01",x"07",x"0d",x"07",x"13",x"07",x"ff",x"09",x"00",x"08",x"01",x"00",
	x"02",x"08",x"02",x"12",x"02",x"00",x"03",x"08",x"03",x"12",x"03",x"00",x"04",x"05",x"04",x"11",
	x"04",x"00",x"05",x"00",x"06",x"05",x"06",x"11",x"06",x"00",x"07",x"06",x"07",x"12",x"07",x"ff",
	x"00",x"00",x"00",x"01",x"00",x"02",x"00",x"03",x"00",x"04",x"00",x"05",x"ff",x"cd",x"0d",x"16",
	x"14",x"32",x"0a",x"64",x"05",x"c8",x"00",x"3e",x"01",x"32",x"44",x"60",x"3a",x"41",x"60",x"dd",
	x"21",x"45",x"60",x"c6",x"0a",x"dd",x"77",x"00",x"dd",x"36",x"01",x"b0",x"18",x"18",x"dd",x"21",
	x"45",x"60",x"21",x"f0",x"0d",x"3e",x"01",x"cd",x"2a",x"14",x"dd",x"7e",x"01",x"d6",x"04",x"fe",
	x"04",x"28",x"16",x"dd",x"77",x"01",x"21",x"f0",x"0d",x"af",x"c3",x"2a",x"14",x"dd",x"21",x"45",
	x"60",x"21",x"f0",x"0d",x"3e",x"01",x"cd",x"2a",x"14",x"af",x"32",x"44",x"60",x"c9",x"dd",x"e5",
	x"e5",x"3e",x"ff",x"32",x"43",x"60",x"3a",x"41",x"60",x"32",x"66",x"60",x"c6",x"28",x"32",x"41",
	x"60",x"cd",x"2e",x"0d",x"cd",x"0d",x"16",x"01",x"0f",x"00",x"3a",x"66",x"60",x"dd",x"be",x"00",
	x"20",x"ef",x"e1",x"dd",x"e1",x"c9",x"0e",x"20",x"5e",x"23",x"56",x"23",x"06",x"0b",x"dd",x"73",
	x"00",x"dd",x"23",x"dd",x"72",x"00",x"dd",x"23",x"10",x"f4",x"0d",x"20",x"eb",x"c9",x"3a",x"29",
	x"60",x"c6",x"03",x"32",x"6a",x"60",x"21",x"af",x"0f",x"22",x"68",x"60",x"3e",x"04",x"32",x"67",
	x"60",x"dd",x"21",x"6b",x"60",x"dd",x"36",x"00",x"05",x"dd",x"23",x"3a",x"6a",x"60",x"dd",x"77",
	x"00",x"dd",x"23",x"3c",x"3c",x"32",x"6a",x"60",x"2a",x"68",x"60",x"7e",x"23",x"22",x"68",x"60",
	x"cd",x"e2",x"0e",x"cd",x"76",x"0e",x"3a",x"67",x"60",x"3d",x"32",x"67",x"60",x"f2",x"a5",x"0e",
	x"c9",x"dd",x"21",x"6b",x"60",x"b7",x"c8",x"c5",x"01",x"c2",x"02",x"dd",x"09",x"3d",x"20",x"fb",
	x"c1",x"c9",x"21",x"ef",x"0e",x"b7",x"c8",x"01",x"40",x"00",x"09",x"3d",x"20",x"fc",x"c9",x"1f",
	x"80",x"3f",x"c0",x"7f",x"e0",x"ff",x"f0",x"de",x"f0",x"de",x"f0",x"de",x"f0",x"ff",x"f0",x"3f",
	x"80",x"30",x"c0",x"60",x"60",x"c0",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1f",
	x"80",x"3f",x"c0",x"7f",x"e0",x"ff",x"f0",x"f7",x"b0",x"f7",x"b0",x"f7",x"b0",x"ff",x"f0",x"1f",
	x"80",x"19",x"80",x"19",x"80",x"19",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c0",
	x"30",x"c0",x"30",x"ff",x"f0",x"86",x"10",x"e7",x"90",x"86",x"10",x"ff",x"f0",x"2f",x"40",x"4f",
	x"20",x"86",x"10",x"40",x"20",x"20",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c0",
	x"30",x"c0",x"30",x"ff",x"f0",x"86",x"10",x"9e",x"70",x"86",x"10",x"ff",x"f0",x"2f",x"40",x"2f",
	x"40",x"26",x"40",x"20",x"40",x"20",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"30",
	x"c0",x"30",x"c0",x"09",x"00",x"0f",x"00",x"1f",x"80",x"3f",x"c0",x"7f",x"e0",x"b0",x"d0",x"9f",
	x"90",x"09",x"00",x"10",x"80",x"09",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c0",
	x"30",x"c0",x"30",x"20",x"40",x"16",x"80",x"1f",x"80",x"3f",x"c0",x"ff",x"f0",x"30",x"c0",x"1f",
	x"80",x"09",x"00",x"10",x"80",x"20",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",
	x"01",x"01",x"00",x"00",x"3a",x"3b",x"60",x"47",x"3a",x"3d",x"60",x"b8",x"30",x"15",x"32",x"3b",
	x"60",x"3a",x"3c",x"60",x"b7",x"20",x"0c",x"3a",x"3b",x"60",x"cd",x"d1",x"0e",x"cd",x"ae",x"10",
	x"cd",x"1a",x"10",x"3a",x"3b",x"60",x"b7",x"20",x"06",x"cd",x"0d",x"16",x"0a",x"fa",x"00",x"cd",
	x"d1",x"0e",x"cd",x"ae",x"10",x"3a",x"3c",x"60",x"b7",x"28",x"1a",x"cd",x"3e",x"10",x"3a",x"3b",
	x"60",x"b7",x"20",x"0c",x"32",x"3c",x"60",x"3a",x"3e",x"60",x"ed",x"44",x"32",x"3e",x"60",x"c9",
	x"3d",x"32",x"3b",x"60",x"c9",x"cd",x"83",x"10",x"3a",x"3b",x"60",x"47",x"3a",x"3d",x"60",x"b8",
	x"28",x"08",x"3a",x"3b",x"60",x"3c",x"32",x"3b",x"60",x"c9",x"3a",x"3e",x"60",x"fe",x"01",x"28",
	x"0c",x"3a",x"39",x"6e",x"b7",x"20",x"12",x"3e",x"01",x"32",x"3c",x"60",x"c9",x"3a",x"39",x"6e",
	x"47",x"3a",x"3a",x"6e",x"80",x"fe",x"20",x"28",x"ee",x"af",x"32",x"3b",x"60",x"c9",x"cd",x"0d",
	x"16",x"08",x"fa",x"00",x"3a",x"38",x"6e",x"fe",x"12",x"d4",x"7e",x"11",x"3a",x"38",x"6e",x"fe",
	x"15",x"28",x"1e",x"47",x"0e",x"00",x"cd",x"f8",x"15",x"cd",x"99",x"0a",x"ed",x"4b",x"37",x"6e",
	x"04",x"dd",x"2a",x"35",x"6e",x"dd",x"71",x"00",x"dd",x"70",x"01",x"cd",x"ae",x"10",x"c3",x"fd",
	x"10",x"3e",x"01",x"32",x"28",x"60",x"cd",x"0d",x"16",x"fa",x"64",x"fa",x"c8",x"fa",x"fa",x"fa",
	x"fa",x"00",x"c9",x"ed",x"4b",x"37",x"6e",x"3a",x"3e",x"60",x"81",x"4f",x"18",x"d3",x"3e",x"04",
	x"32",x"3b",x"60",x"cd",x"d1",x"0e",x"cd",x"ae",x"10",x"cd",x"fd",x"10",x"cd",x"0d",x"16",x"19",
	x"f0",x"64",x"78",x"19",x"f0",x"00",x"3a",x"3b",x"60",x"3d",x"f2",x"90",x"10",x"c9",x"dd",x"22",
	x"35",x"6e",x"dd",x"4e",x"00",x"dd",x"46",x"01",x"ed",x"43",x"37",x"6e",x"3a",x"3f",x"60",x"3c",
	x"cb",x"27",x"4f",x"06",x"00",x"dd",x"09",x"3a",x"37",x"6e",x"1f",x"30",x"05",x"01",x"60",x"01",
	x"dd",x"09",x"dd",x"22",x"3c",x"6e",x"3a",x"37",x"6e",x"47",x"3a",x"3f",x"60",x"cb",x"27",x"80",
	x"32",x"39",x"6e",x"3a",x"3f",x"60",x"47",x"3a",x"40",x"60",x"90",x"cb",x"27",x"32",x"3a",x"6e",
	x"47",x"3a",x"39",x"6e",x"80",x"d6",x"20",x"ed",x"44",x"32",x"3b",x"6e",x"c9",x"cd",x"66",x"11",
	x"ed",x"4b",x"37",x"6e",x"cd",x"0c",x"11",x"ed",x"4b",x"37",x"6e",x"04",x"3e",x"08",x"32",x"40",
	x"6e",x"0e",x"00",x"cd",x"f8",x"15",x"ed",x"53",x"3e",x"6e",x"cd",x"38",x"11",x"2a",x"3c",x"6e",
	x"01",x"16",x"00",x"09",x"22",x"3c",x"6e",x"2a",x"3e",x"6e",x"24",x"22",x"3e",x"6e",x"3a",x"40",
	x"6e",x"3d",x"32",x"40",x"6e",x"20",x"e3",x"c9",x"ed",x"5b",x"3e",x"6e",x"3a",x"39",x"6e",x"cd",
	x"50",x"11",x"2a",x"3c",x"6e",x"ed",x"4b",x"3a",x"6e",x"06",x"00",x"ed",x"b0",x"3a",x"3b",x"6e",
	x"b7",x"c8",x"47",x"af",x"12",x"13",x"10",x"fc",x"c9",x"cd",x"41",x"13",x"3e",x"f8",x"a6",x"b3",
	x"77",x"23",x"15",x"20",x"f7",x"c9",x"ed",x"4b",x"37",x"6e",x"0e",x"00",x"21",x"3b",x"05",x"3a",
	x"3b",x"60",x"85",x"6f",x"30",x"01",x"24",x"7e",x"5f",x"16",x"40",x"c3",x"59",x"11",x"3a",x"25",
	x"60",x"b7",x"c8",x"11",x"80",x"50",x"cd",x"99",x"0a",x"11",x"a0",x"50",x"cd",x"99",x"0a",x"11",
	x"c0",x"50",x"cd",x"99",x"0a",x"af",x"32",x"25",x"60",x"cd",x"0d",x"16",x"c8",x"0a",x"0a",x"c8",
	x"c8",x"0a",x"0a",x"c8",x"c8",x"0a",x"32",x"fa",x"00",x"c9",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"03",x"0f",x"1f",x"3f",x"7f",x"7f",x"ff",x"ff",x"c0",x"f0",x"f8",x"fc",x"fe",x"fe",
	x"ff",x"ff",x"fc",x"f0",x"e0",x"c0",x"80",x"80",x"00",x"00",x"3f",x"0f",x"07",x"03",x"01",x"01",
	x"00",x"00",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"00",x"00",x"31",x"30",x"30",x"32",x"00",x"30",
	x"30",x"30",x"30",x"00",x"35",x"33",x"34",x"35",x"00",x"3a",x"25",x"60",x"b7",x"c0",x"2a",x"1a",
	x"60",x"e5",x"21",x"2a",x"10",x"22",x"1a",x"60",x"3e",x"03",x"32",x"41",x"6e",x"01",x"05",x"14",
	x"21",x"da",x"11",x"c5",x"3e",x"03",x"32",x"42",x"6e",x"cd",x"91",x"15",x"0d",x"0d",x"0d",x"0d",
	x"04",x"3a",x"42",x"6e",x"3d",x"32",x"42",x"6e",x"20",x"ef",x"c1",x"79",x"c6",x"09",x"4f",x"3a",
	x"41",x"6e",x"3d",x"32",x"41",x"6e",x"20",x"d8",x"e1",x"22",x"1a",x"60",x"3e",x"01",x"32",x"25",
	x"60",x"c9",x"fe",x"00",x"ff",x"00",x"01",x"00",x"02",x"00",x"ff",x"ff",x"01",x"ff",x"ff",x"01",
	x"01",x"01",x"3a",x"25",x"60",x"b7",x"c8",x"ed",x"43",x"43",x"6e",x"78",x"fe",x"a2",x"38",x"5b",
	x"fe",x"b8",x"30",x"57",x"cd",x"55",x"14",x"c8",x"cd",x"b6",x"18",x"dd",x"21",x"32",x"12",x"3e",
	x"08",x"32",x"41",x"6e",x"3a",x"43",x"6e",x"dd",x"86",x"00",x"4f",x"3a",x"44",x"6e",x"dd",x"86",
	x"01",x"47",x"dd",x"23",x"dd",x"23",x"3a",x"a4",x"6e",x"17",x"32",x"a4",x"6e",x"dc",x"48",x"14",
	x"3a",x"41",x"6e",x"3d",x"32",x"41",x"6e",x"20",x"db",x"ed",x"4b",x"43",x"6e",x"cd",x"48",x"14",
	x"ed",x"4b",x"43",x"6e",x"04",x"cd",x"48",x"14",x"ed",x"4b",x"43",x"6e",x"05",x"cd",x"48",x"14",
	x"cd",x"0d",x"16",x"04",x"14",x"04",x"1e",x"00",x"f6",x"01",x"c9",x"af",x"c9",x"21",x"00",x"40",
	x"0e",x"18",x"af",x"47",x"77",x"23",x"10",x"fc",x"0d",x"20",x"f9",x"c9",x"10",x"27",x"e8",x"03",
	x"64",x"00",x"0a",x"00",x"01",x"00",x"dd",x"21",x"45",x"6e",x"06",x"05",x"ed",x"73",x"4a",x"6e",
	x"31",x"bc",x"12",x"d1",x"f6",x"ff",x"ed",x"52",x"3c",x"30",x"fb",x"19",x"dd",x"77",x"00",x"dd",
	x"23",x"10",x"f0",x"dd",x"21",x"45",x"6e",x"ed",x"7b",x"4a",x"6e",x"c9",x"11",x"01",x"01",x"22",
	x"4c",x"6e",x"79",x"95",x"d2",x"fb",x"12",x"1e",x"ff",x"ed",x"44",x"4f",x"78",x"94",x"d2",x"05",
	x"13",x"16",x"ff",x"ed",x"44",x"47",x"79",x"b8",x"30",x"06",x"69",x"d5",x"af",x"5f",x"18",x"07",
	x"b1",x"c8",x"68",x"41",x"d5",x"16",x"00",x"60",x"78",x"1f",x"85",x"38",x"03",x"bc",x"38",x"07",
	x"94",x"4f",x"d9",x"c1",x"c5",x"18",x"04",x"4f",x"d5",x"d9",x"c1",x"2a",x"4c",x"6e",x"78",x"84",
	x"47",x"79",x"85",x"4f",x"ed",x"43",x"4c",x"6e",x"cd",x"5e",x"13",x"d9",x"79",x"10",x"db",x"d1",
	x"c9",x"78",x"f6",x"c0",x"6f",x"26",x"02",x"29",x"29",x"29",x"29",x"29",x"79",x"85",x"6f",x"d0",
	x"24",x"c9",x"cd",x"f8",x"15",x"06",x"08",x"7e",x"23",x"12",x"14",x"10",x"fa",x"c9",x"2a",x"4e",
	x"6e",x"e9",x"42",x"14",x"48",x"14",x"4f",x"14",x"55",x"14",x"e5",x"c5",x"e6",x"03",x"6f",x"26",
	x"00",x"29",x"01",x"62",x"13",x"09",x"01",x"4e",x"6e",x"7e",x"02",x"23",x"03",x"7e",x"02",x"c1",
	x"e1",x"c9",x"a7",x"f2",x"8f",x"13",x"21",x"00",x"00",x"b7",x"ed",x"52",x"eb",x"ed",x"44",x"4b",
	x"5a",x"16",x"00",x"47",x"cb",x"7b",x"28",x"01",x"15",x"62",x"cb",x"21",x"cb",x"13",x"cb",x"12",
	x"79",x"cb",x"17",x"7b",x"6a",x"cb",x"17",x"cb",x"15",x"cb",x"14",x"81",x"4f",x"ed",x"5a",x"eb",
	x"21",x"00",x"00",x"78",x"06",x"07",x"cb",x"1f",x"30",x"08",x"19",x"cb",x"21",x"30",x"05",x"23",
	x"18",x"02",x"cb",x"21",x"cb",x"13",x"cb",x"12",x"10",x"ec",x"c9",x"21",x"da",x"13",x"cb",x"27",
	x"cb",x"27",x"cb",x"27",x"85",x"6f",x"30",x"01",x"24",x"c9",x"7e",x"7e",x"66",x"66",x"66",x"66",
	x"7e",x"7e",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"7e",x"7e",x"06",x"7e",x"7e",x"60",
	x"7e",x"7e",x"7e",x"7e",x"06",x"7e",x"7e",x"06",x"7e",x"7e",x"60",x"60",x"6c",x"6c",x"7e",x"7e",
	x"0c",x"0c",x"7e",x"7e",x"60",x"7e",x"7e",x"06",x"7e",x"7e",x"7e",x"7e",x"60",x"7e",x"7e",x"66",
	x"7e",x"7e",x"7e",x"7e",x"06",x"06",x"06",x"06",x"06",x"06",x"7e",x"7e",x"66",x"7e",x"7e",x"66",
	x"7e",x"7e",x"7e",x"7e",x"66",x"7e",x"7e",x"06",x"7e",x"7e",x"cd",x"6a",x"13",x"7e",x"23",x"b7",
	x"f8",x"dd",x"86",x"00",x"4f",x"7e",x"23",x"dd",x"86",x"01",x"47",x"e5",x"cd",x"5e",x"13",x"e1",
	x"18",x"eb",x"cd",x"62",x"15",x"b6",x"77",x"c9",x"cd",x"62",x"15",x"2f",x"a6",x"77",x"c9",x"cd",
	x"62",x"15",x"ae",x"77",x"c9",x"cd",x"62",x"15",x"a6",x"c9",x"80",x"40",x"20",x"10",x"08",x"04",
	x"02",x"01",x"00",x"08",x"10",x"18",x"20",x"28",x"30",x"38",x"01",x"09",x"11",x"19",x"21",x"29",
	x"31",x"39",x"02",x"0a",x"12",x"1a",x"22",x"2a",x"32",x"3a",x"03",x"0b",x"13",x"1b",x"23",x"2b",
	x"33",x"3b",x"04",x"0c",x"14",x"1c",x"24",x"2c",x"34",x"3c",x"05",x"0d",x"15",x"1d",x"25",x"2d",
	x"35",x"3d",x"06",x"0e",x"16",x"1e",x"26",x"2e",x"36",x"3e",x"07",x"0f",x"17",x"1f",x"27",x"2f",
	x"37",x"3f",x"40",x"48",x"50",x"58",x"60",x"68",x"70",x"78",x"41",x"49",x"51",x"59",x"61",x"69",
	x"71",x"79",x"42",x"4a",x"52",x"5a",x"62",x"6a",x"72",x"7a",x"43",x"4b",x"53",x"5b",x"63",x"6b",
	x"73",x"7b",x"44",x"4c",x"54",x"5c",x"64",x"6c",x"74",x"7c",x"45",x"4d",x"55",x"5d",x"65",x"6d",
	x"75",x"7d",x"46",x"4e",x"56",x"5e",x"66",x"6e",x"76",x"7e",x"47",x"4f",x"57",x"5f",x"67",x"6f",
	x"77",x"7f",x"80",x"88",x"90",x"98",x"a0",x"a8",x"b0",x"b8",x"81",x"89",x"91",x"99",x"a1",x"a9",
	x"b1",x"b9",x"82",x"8a",x"92",x"9a",x"a2",x"aa",x"b2",x"ba",x"83",x"8b",x"93",x"9b",x"a3",x"ab",
	x"b3",x"bb",x"84",x"8c",x"94",x"9c",x"a4",x"ac",x"b4",x"bc",x"85",x"8d",x"95",x"9d",x"a5",x"ad",
	x"b5",x"bd",x"86",x"8e",x"96",x"9e",x"a6",x"ae",x"b6",x"be",x"87",x"8f",x"97",x"9f",x"a7",x"af",
	x"b7",x"bf",x"00",x"08",x"10",x"18",x"20",x"28",x"30",x"38",x"01",x"09",x"11",x"19",x"21",x"29",
	x"31",x"39",x"02",x"0a",x"12",x"1a",x"22",x"2a",x"32",x"3a",x"03",x"0b",x"13",x"1b",x"23",x"2b",
	x"33",x"3b",x"84",x"8c",x"94",x"9c",x"a4",x"ac",x"b4",x"bc",x"85",x"8d",x"95",x"9d",x"a5",x"ad",
	x"b5",x"bd",x"86",x"8e",x"96",x"9e",x"a6",x"ae",x"b6",x"be",x"87",x"8f",x"97",x"9f",x"a7",x"af",
	x"b7",x"bf",x"21",x"62",x"14",x"58",x"16",x"00",x"19",x"66",x"69",x"a7",x"cb",x"1c",x"cb",x"1d",
	x"37",x"cb",x"1c",x"cb",x"1d",x"a7",x"cb",x"1c",x"cb",x"1d",x"eb",x"21",x"5a",x"14",x"79",x"e6",
	x"07",x"4f",x"06",x"00",x"09",x"7e",x"eb",x"c9",x"e1",x"cd",x"8d",x"15",x"e9",x"4e",x"23",x"46",
	x"23",x"7e",x"23",x"b7",x"c8",x"fe",x"01",x"28",x"f4",x"c5",x"e5",x"cd",x"eb",x"18",x"cd",x"52",
	x"13",x"e1",x"c1",x"cd",x"a8",x"15",x"18",x"e9",x"0c",x"79",x"fe",x"20",x"c0",x"0e",x"00",x"04",
	x"78",x"fe",x"18",x"c0",x"06",x"00",x"c9",x"e1",x"ed",x"73",x"50",x"6e",x"31",x"85",x"6e",x"e5",
	x"fd",x"22",x"86",x"6e",x"d9",x"22",x"88",x"6e",x"ed",x"53",x"8a",x"6e",x"ed",x"43",x"8c",x"6e",
	x"d9",x"c9",x"ed",x"73",x"52",x"6e",x"ed",x"7b",x"50",x"6e",x"d9",x"2a",x"88",x"6e",x"ed",x"5b",
	x"8a",x"6e",x"ed",x"4b",x"8c",x"6e",x"d9",x"fd",x"2a",x"86",x"6e",x"fb",x"c9",x"ed",x"73",x"50",
	x"6e",x"ed",x"7b",x"52",x"6e",x"c3",x"c4",x"15",x"50",x"af",x"cb",x"18",x"1f",x"cb",x"18",x"1f",
	x"cb",x"18",x"1f",x"b1",x"5f",x"42",x"3e",x"18",x"a2",x"f6",x"40",x"57",x"c9",x"ed",x"53",x"8e",
	x"6e",x"d1",x"c5",x"f5",x"e5",x"3a",x"48",x"5c",x"e6",x"38",x"0f",x"0f",x"0f",x"f6",x"08",x"32",
	x"90",x"6e",x"1a",x"13",x"b7",x"28",x"09",x"6f",x"1a",x"13",x"67",x"cd",x"39",x"16",x"18",x"f2",
	x"e1",x"f1",x"c1",x"d5",x"ed",x"5b",x"8e",x"6e",x"c9",x"cd",x"40",x"16",x"2d",x"20",x"fa",x"c9",
	x"3a",x"90",x"6e",x"cd",x"4a",x"16",x"06",x"04",x"10",x"fe",x"44",x"00",x"00",x"00",x"10",x"fb",
	x"ee",x"10",x"d3",x"fe",x"c9",x"00",x"01",x"02",x"02",x"03",x"04",x"05",x"05",x"06",x"07",x"08",
	x"09",x"09",x"0a",x"0b",x"0c",x"0c",x"0d",x"0e",x"0f",x"10",x"10",x"11",x"12",x"13",x"13",x"14",
	x"15",x"16",x"17",x"17",x"18",x"19",x"1a",x"1a",x"1b",x"1c",x"1d",x"1d",x"1e",x"1f",x"20",x"20",
	x"21",x"22",x"23",x"24",x"24",x"25",x"26",x"27",x"27",x"28",x"29",x"29",x"2a",x"2b",x"2c",x"2c",
	x"2d",x"2e",x"2f",x"2f",x"30",x"31",x"32",x"32",x"33",x"34",x"34",x"35",x"36",x"36",x"37",x"38",
	x"39",x"39",x"3a",x"3b",x"3b",x"3c",x"3d",x"3d",x"3e",x"3f",x"40",x"40",x"41",x"42",x"42",x"43",
	x"44",x"44",x"45",x"45",x"46",x"47",x"47",x"48",x"49",x"49",x"4a",x"4b",x"4b",x"4c",x"4d",x"4d",
	x"4e",x"4e",x"4f",x"50",x"50",x"51",x"51",x"52",x"53",x"53",x"54",x"54",x"55",x"56",x"56",x"57",
	x"57",x"58",x"58",x"59",x"5a",x"5a",x"5b",x"5b",x"5c",x"5c",x"5d",x"5d",x"5e",x"5e",x"5f",x"5f",
	x"60",x"60",x"61",x"61",x"62",x"62",x"63",x"63",x"64",x"64",x"65",x"65",x"66",x"66",x"67",x"67",
	x"68",x"68",x"69",x"69",x"69",x"6a",x"6a",x"6b",x"6b",x"6c",x"6c",x"6c",x"6d",x"6d",x"6e",x"6e",
	x"6e",x"6f",x"6f",x"70",x"70",x"70",x"71",x"71",x"71",x"72",x"72",x"72",x"73",x"73",x"73",x"74",
	x"74",x"74",x"75",x"75",x"75",x"76",x"76",x"76",x"76",x"77",x"77",x"77",x"78",x"78",x"78",x"78",
	x"79",x"79",x"79",x"79",x"79",x"7a",x"7a",x"7a",x"7a",x"7b",x"7b",x"7b",x"7b",x"7b",x"7c",x"7c",
	x"7c",x"7c",x"7c",x"7c",x"7d",x"7d",x"7d",x"7d",x"7d",x"7d",x"7d",x"7d",x"7e",x"7e",x"7e",x"7e",
	x"7e",x"7e",x"7e",x"7e",x"7e",x"7e",x"7f",x"7f",x"7f",x"7f",x"7f",x"7f",x"7f",x"7f",x"7f",x"7f",
	x"7f",x"7f",x"7f",x"7f",x"7f",x"01",x"fc",x"03",x"cb",x"7c",x"28",x"04",x"09",x"30",x"fd",x"c9",
	x"b7",x"ed",x"42",x"30",x"fc",x"09",x"c9",x"cd",x"55",x"17",x"01",x"ff",x"00",x"b7",x"ed",x"42",
	x"30",x"03",x"09",x"18",x"21",x"ed",x"42",x"30",x"08",x"7d",x"ed",x"44",x"6f",x"26",x"00",x"18",
	x"15",x"ed",x"42",x"38",x"0a",x"ed",x"42",x"7d",x"ed",x"44",x"6f",x"26",x"00",x"18",x"01",x"09",
	x"cd",x"96",x"17",x"ed",x"44",x"c9",x"01",x"55",x"16",x"09",x"7e",x"c9",x"24",x"2b",x"c3",x"67",
	x"17",x"2a",x"a2",x"6e",x"7e",x"23",x"22",x"91",x"6e",x"6f",x"3c",x"c8",x"26",x"00",x"29",x"29",
	x"29",x"ed",x"4b",x"1a",x"60",x"09",x"3e",x"08",x"32",x"95",x"6e",x"3a",x"9e",x"6e",x"32",x"9a",
	x"6e",x"3a",x"9d",x"6e",x"32",x"99",x"6e",x"3e",x"09",x"32",x"96",x"6e",x"7e",x"23",x"22",x"93",
	x"6e",x"07",x"32",x"97",x"6e",x"3a",x"96",x"6e",x"3d",x"20",x"32",x"3a",x"95",x"6e",x"3d",x"20",
	x"18",x"3a",x"a1",x"6e",x"47",x"3a",x"9f",x"6e",x"4f",x"3a",x"9d",x"6e",x"81",x"05",x"20",x"fc",
	x"32",x"9d",x"6e",x"2a",x"91",x"6e",x"c3",x"a4",x"17",x"32",x"95",x"6e",x"3a",x"a0",x"6e",x"47",
	x"3a",x"9a",x"6e",x"80",x"32",x"9a",x"6e",x"2a",x"93",x"6e",x"c3",x"c1",x"17",x"32",x"96",x"6e",
	x"3a",x"9f",x"6e",x"47",x"3a",x"9a",x"6e",x"32",x"98",x"6e",x"3a",x"a0",x"6e",x"4f",x"c5",x"cd",
	x"45",x"18",x"c1",x"3a",x"98",x"6e",x"3c",x"32",x"98",x"6e",x"0d",x"20",x"f1",x"3a",x"99",x"6e",
	x"3c",x"32",x"99",x"6e",x"05",x"20",x"dd",x"3a",x"97",x"6e",x"c3",x"d1",x"17",x"80",x"40",x"20",
	x"10",x"08",x"04",x"02",x"01",x"3a",x"9c",x"6e",x"ee",x"ff",x"47",x"3a",x"9b",x"6e",x"a0",x"47",
	x"3a",x"99",x"6e",x"e6",x"f8",x"6f",x"3a",x"98",x"6e",x"fe",x"c0",x"d0",x"1f",x"1f",x"1f",x"e6",
	x"1f",x"67",x"cb",x"1c",x"cb",x"1d",x"cb",x"1c",x"cb",x"1d",x"cb",x"1c",x"cb",x"1d",x"3e",x"58",
	x"b4",x"67",x"3a",x"9c",x"6e",x"a6",x"b0",x"77",x"3a",x"98",x"6e",x"47",x"e6",x"07",x"f6",x"40",
	x"67",x"78",x"1f",x"1f",x"1f",x"e6",x"18",x"b4",x"67",x"78",x"17",x"17",x"e6",x"e0",x"6f",x"3a",
	x"99",x"6e",x"47",x"1f",x"1f",x"1f",x"e6",x"1f",x"b5",x"6f",x"eb",x"21",x"3d",x"18",x"78",x"e6",
	x"07",x"4f",x"06",x"00",x"09",x"46",x"1a",x"21",x"97",x"6e",x"cb",x"46",x"28",x"03",x"b0",x"12",
	x"c9",x"2f",x"b0",x"2f",x"12",x"c9",x"2a",x"a6",x"6e",x"cb",x"15",x"cb",x"14",x"cb",x"15",x"cb",
	x"14",x"4c",x"3a",x"a4",x"6e",x"17",x"47",x"ed",x"5b",x"a5",x"6e",x"cb",x"13",x"cb",x"12",x"cb",
	x"ba",x"2a",x"a4",x"6e",x"09",x"22",x"a4",x"6e",x"2a",x"a6",x"6e",x"ed",x"5a",x"cb",x"bc",x"22",
	x"a6",x"6e",x"f0",x"21",x"a4",x"6e",x"34",x"c0",x"34",x"18",x"fb",x"c5",x"6f",x"26",x"00",x"29",
	x"29",x"29",x"ed",x"4b",x"1a",x"60",x"09",x"c1",x"c9",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
	x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",


	others => x"07"
);

signal ReadAddress: std_logic_vector(Address'range);
signal DualReadAddress: std_logic_vector(DualAddress'range);

attribute syn_ramstyle: string;
attribute syn_ramstyle of RAM: signal is "block_ram";

begin

	process (Clock)
	begin
		if rising_edge(Clock) then
			if Enable = '1' and WriteEnable = '1' then
				RAM(conv_integer(Address)) <= DataIn;
			end if;

			if Enable = '1' then
				ReadAddress <= Address;
			end if;
			if DualEnable = '1' then
				DualReadAddress <= DualAddress;
			end if;
		end if;
	end process;

	DataOut <= RAM(conv_integer(ReadAddress));
	DualDataOut <= RAM(conv_integer(DualReadAddress));

end behavioral;
